** Generated for: hspiceD
** Generated on: Jan 26 16:01:37 2024
** Design library name: ising
** Design cell name: ising_50x50
** Design view name: schematic

** Library name: ising
** Cell name: unit_coupling_tile
** View name: schematic
.subckt unit_coupling_tile d2u_in d2u_out l2r_in l2r_out r2l_in r2l_out u2d_in u2d_out vdd vss
.ends unit_coupling_tile
** End of subcircuit definition.

** Library name: ising
** Cell name: short_tile
** View name: schematic
.subckt short_tile d2u_in d2u_out l2r_in l2r_out r2l_in r2l_out u2d_in u2d_out vdd vss
.ends short_tile
** End of subcircuit definition.

** Library name: ising
** Cell name: enable_tile
** View name: schematic
.subckt enable_tile vdd vss enable in_ out_
.ends enable_tile
** End of subcircuit definition.

** Library name: ising
** Cell name: ising_50x50
** View name: schematic
xi2499 net10342 net10175 net10306 net53 net53 net10303 net10174 net10341 vdd vss unit_coupling_tile
xi2498 net10305 net10173 net10302 net10306 net10303 net10299 net10172 net10304 vdd vss unit_coupling_tile
xi2497 net10301 net10101 net10312 net10302 net10299 net10309 net10100 net10300 vdd vss unit_coupling_tile
xi2496 net10311 net10097 net10313 net10312 net10309 net10307 net10096 net10310 vdd vss unit_coupling_tile
xi2495 net10320 net10107 net10317 net10313 net10307 net10314 net10106 net10308 vdd vss unit_coupling_tile
xi2494 net10316 net10116 net10318 net10317 net10314 net10319 net10104 net10315 vdd vss unit_coupling_tile
xi2493 net10325 net10112 net10326 net10318 net10319 net10321 net10111 net10324 vdd vss unit_coupling_tile
xi2492 net10323 net10121 net10330 net10326 net10321 net10327 net10120 net10322 vdd vss unit_coupling_tile
xi2491 net10329 net10119 net10331 net10330 net10327 net10332 net10118 net10328 vdd vss unit_coupling_tile
xi2490 net10338 net10125 net10336 net10331 net10332 net10333 net10124 net10337 vdd vss unit_coupling_tile
xi2489 net10335 net10134 net10265 net10336 net10333 net10339 net10133 net10334 vdd vss unit_coupling_tile
xi2488 net10264 net10131 net10261 net10265 net10339 net10258 net10130 net10340 vdd vss unit_coupling_tile
xi2487 net10260 net10060 net10262 net10261 net10258 net10263 net10136 net10259 vdd vss unit_coupling_tile
xi2486 net10270 net10056 net10271 net10262 net10263 net10266 net10055 net10269 vdd vss unit_coupling_tile
xi2485 net10268 net10066 net10275 net10271 net10266 net10272 net10065 net10267 vdd vss unit_coupling_tile
xi2484 net10274 net10064 net10276 net10275 net10272 net10277 net10063 net10273 vdd vss unit_coupling_tile
xi2483 net10283 net10070 net10281 net10276 net10277 net10278 net10069 net10282 vdd vss unit_coupling_tile
xi2482 net10280 net10079 net10289 net10281 net10278 net10286 net10078 net10279 vdd vss unit_coupling_tile
xi2481 net10288 net10076 net10290 net10289 net10286 net10284 net10075 net10287 vdd vss unit_coupling_tile
xi2480 net10296 net10084 net10294 net10290 net10284 net10291 net10083 net10285 vdd vss unit_coupling_tile
xi2479 net10293 net10092 net10223 net10294 net10291 net10295 net10081 net10292 vdd vss unit_coupling_tile
xi2478 net10298 net10089 net10220 net10223 net10295 net10217 net10088 net10297 vdd vss unit_coupling_tile
xi2477 net10219 net10094 net10221 net10220 net10217 net10222 net10093 net10218 vdd vss unit_coupling_tile
xi2476 net10229 net10015 net10227 net10221 net10222 net10224 net10014 net10228 vdd vss unit_coupling_tile
xi2475 net10226 net10025 net10235 net10227 net10224 net10232 net10024 net10225 vdd vss unit_coupling_tile
xi2474 net10234 net10022 net10236 net10235 net10232 net10230 net10021 net10233 vdd vss unit_coupling_tile
xi2473 net10243 net10030 net10240 net10236 net10230 net10237 net10029 net10231 vdd vss unit_coupling_tile
xi2472 net10239 net10039 net10241 net10240 net10237 net10242 net10027 net10238 vdd vss unit_coupling_tile
xi2471 net10248 net10035 net10249 net10241 net10242 net10244 net10034 net10247 vdd vss unit_coupling_tile
xi2470 net10246 net10044 net10253 net10249 net10244 net10250 net10043 net10245 vdd vss unit_coupling_tile
xi2469 net10252 net10042 net10254 net10253 net10250 net10255 net10041 net10251 vdd vss unit_coupling_tile
xi2468 net10257 net10048 net10182 net10254 net10255 net10179 net10047 net10256 vdd vss unit_coupling_tile
xi2467 net10181 net10053 net10183 net10182 net10179 net10177 net10052 net10180 vdd vss unit_coupling_tile
xi2466 net10190 net9977 net10187 net10183 net10177 net10184 net9976 net10178 vdd vss unit_coupling_tile
xi2465 net10186 net9986 net10188 net10187 net10184 net10189 net9974 net10185 vdd vss unit_coupling_tile
xi2464 net10195 net9982 net10196 net10188 net10189 net10191 net9981 net10194 vdd vss unit_coupling_tile
xi2463 net10193 net9991 net10200 net10196 net10191 net10197 net9990 net10192 vdd vss unit_coupling_tile
xi2462 net10199 net9989 net10201 net10200 net10197 net10202 net9988 net10198 vdd vss unit_coupling_tile
xi2461 net10208 net9995 net10206 net10201 net10202 net10203 net9994 net10207 vdd vss unit_coupling_tile
xi2460 net10205 net10004 net10214 net10206 net10203 net10211 net10003 net10204 vdd vss unit_coupling_tile
xi2459 net10213 net10001 net10215 net10214 net10211 net10209 net10000 net10212 vdd vss unit_coupling_tile
xi2458 net10216 net10009 net10143 net10215 net10209 net10140 net10008 net10210 vdd vss unit_coupling_tile
xi2457 net10142 net10012 net10144 net10143 net10140 net10137 net10006 net10141 vdd vss unit_coupling_tile
xi2456 net10139 net9938 net10148 net10144 net10137 net10145 net9937 net10138 vdd vss unit_coupling_tile
xi2455 net10147 net9935 net10149 net10148 net10145 net10150 net9934 net10146 vdd vss unit_coupling_tile
xi2454 net10156 net9943 net10154 net10149 net10150 net10151 net9942 net10155 vdd vss unit_coupling_tile
xi2453 net10153 net9952 net10162 net10154 net10151 net10159 net9951 net10152 vdd vss unit_coupling_tile
xi2452 net10161 net9949 net10163 net10162 net10159 net10157 net9948 net10160 vdd vss unit_coupling_tile
xi2451 net10164 net9958 net10165 net10163 net10157 net10166 net9957 net10158 vdd vss unit_coupling_tile
xi2449 net10175 net9961 net10176 net54 net54 net10171 net9960 net10174 vdd vss unit_coupling_tile
xi2448 net10173 net9971 net10102 net10176 net10171 net10099 net9970 net10172 vdd vss unit_coupling_tile
xi2447 net10101 net9969 net10098 net10102 net10099 net10095 net9968 net10100 vdd vss unit_coupling_tile
xi2446 net10097 net9897 net10108 net10098 net10095 net10105 net9896 net10096 vdd vss unit_coupling_tile
xi2445 net10107 net9893 net10109 net10108 net10105 net10103 net9892 net10106 vdd vss unit_coupling_tile
xi2444 net10116 net9903 net10113 net10109 net10103 net10110 net9902 net10104 vdd vss unit_coupling_tile
xi2443 net10112 net9912 net10114 net10113 net10110 net10115 net9900 net10111 vdd vss unit_coupling_tile
xi2442 net10121 net9908 net10122 net10114 net10115 net10117 net9907 net10120 vdd vss unit_coupling_tile
xi2441 net10119 net9917 net10126 net10122 net10117 net10123 net9916 net10118 vdd vss unit_coupling_tile
xi2440 net10125 net9915 net10127 net10126 net10123 net10128 net9914 net10124 vdd vss unit_coupling_tile
xi2439 net10134 net9921 net10132 net10127 net10128 net10129 net9920 net10133 vdd vss unit_coupling_tile
xi2438 net10131 net9930 net10061 net10132 net10129 net10135 net9929 net10130 vdd vss unit_coupling_tile
xi2437 net10060 net9927 net10057 net10061 net10135 net10054 net9926 net10136 vdd vss unit_coupling_tile
xi2436 net10056 net9856 net10058 net10057 net10054 net10059 net9932 net10055 vdd vss unit_coupling_tile
xi2435 net10066 net9852 net10067 net10058 net10059 net10062 net9851 net10065 vdd vss unit_coupling_tile
xi2434 net10064 net9862 net10071 net10067 net10062 net10068 net9861 net10063 vdd vss unit_coupling_tile
xi2433 net10070 net9860 net10072 net10071 net10068 net10073 net9859 net10069 vdd vss unit_coupling_tile
xi2432 net10079 net9866 net10077 net10072 net10073 net10074 net9865 net10078 vdd vss unit_coupling_tile
xi2431 net10076 net9875 net10085 net10077 net10074 net10082 net9874 net10075 vdd vss unit_coupling_tile
xi2430 net10084 net9872 net10086 net10085 net10082 net10080 net9871 net10083 vdd vss unit_coupling_tile
xi2429 net10092 net9880 net10090 net10086 net10080 net10087 net9879 net10081 vdd vss unit_coupling_tile
xi2428 net10089 net9888 net10019 net10090 net10087 net10091 net9877 net10088 vdd vss unit_coupling_tile
xi2427 net10094 net9885 net10016 net10019 net10091 net10013 net9884 net10093 vdd vss unit_coupling_tile
xi2426 net10015 net9890 net10017 net10016 net10013 net10018 net9889 net10014 vdd vss unit_coupling_tile
xi2425 net10025 net9811 net10023 net10017 net10018 net10020 net9810 net10024 vdd vss unit_coupling_tile
xi2424 net10022 net9821 net10031 net10023 net10020 net10028 net9820 net10021 vdd vss unit_coupling_tile
xi2423 net10030 net9818 net10032 net10031 net10028 net10026 net9817 net10029 vdd vss unit_coupling_tile
xi2422 net10039 net9826 net10036 net10032 net10026 net10033 net9825 net10027 vdd vss unit_coupling_tile
xi2421 net10035 net9835 net10037 net10036 net10033 net10038 net9823 net10034 vdd vss unit_coupling_tile
xi2420 net10044 net9831 net10045 net10037 net10038 net10040 net9830 net10043 vdd vss unit_coupling_tile
xi2419 net10042 net9840 net10049 net10045 net10040 net10046 net9839 net10041 vdd vss unit_coupling_tile
xi2418 net10048 net9838 net10050 net10049 net10046 net10051 net9837 net10047 vdd vss unit_coupling_tile
xi2417 net10053 net9844 net9978 net10050 net10051 net9975 net9843 net10052 vdd vss unit_coupling_tile
xi2416 net9977 net9849 net9979 net9978 net9975 net9973 net9848 net9976 vdd vss unit_coupling_tile
xi2415 net9986 net9773 net9983 net9979 net9973 net9980 net9772 net9974 vdd vss unit_coupling_tile
xi2414 net9982 net9782 net9984 net9983 net9980 net9985 net9770 net9981 vdd vss unit_coupling_tile
xi2413 net9991 net9778 net9992 net9984 net9985 net9987 net9777 net9990 vdd vss unit_coupling_tile
xi2412 net9989 net9787 net9996 net9992 net9987 net9993 net9786 net9988 vdd vss unit_coupling_tile
xi2411 net9995 net9785 net9997 net9996 net9993 net9998 net9784 net9994 vdd vss unit_coupling_tile
xi2410 net10004 net9791 net10002 net9997 net9998 net9999 net9790 net10003 vdd vss unit_coupling_tile
xi2409 net10001 net9800 net10010 net10002 net9999 net10007 net9799 net10000 vdd vss unit_coupling_tile
xi2408 net10009 net9797 net10011 net10010 net10007 net10005 net9796 net10008 vdd vss unit_coupling_tile
xi2407 net10012 net9805 net9939 net10011 net10005 net9936 net9804 net10006 vdd vss unit_coupling_tile
xi2406 net9938 net9808 net9940 net9939 net9936 net9933 net9802 net9937 vdd vss unit_coupling_tile
xi2405 net9935 net9734 net9944 net9940 net9933 net9941 net9733 net9934 vdd vss unit_coupling_tile
xi2404 net9943 net9731 net9945 net9944 net9941 net9946 net9730 net9942 vdd vss unit_coupling_tile
xi2403 net9952 net9739 net9950 net9945 net9946 net9947 net9738 net9951 vdd vss unit_coupling_tile
xi2402 net9949 net9748 net9955 net9950 net9947 net9956 net9747 net9948 vdd vss unit_coupling_tile
xi2400 net9964 net9752 net9965 net9959 net9953 net9966 net9751 net9954 vdd vss unit_coupling_tile
xi2399 net9961 net9762 net9962 net55 net55 net9963 net9749 net9960 vdd vss unit_coupling_tile
xi2398 net9971 net9758 net9972 net9962 net9963 net9967 net9757 net9970 vdd vss unit_coupling_tile
xi2397 net9969 net9767 net9898 net9972 net9967 net9895 net9766 net9968 vdd vss unit_coupling_tile
xi2396 net9897 net9765 net9894 net9898 net9895 net9891 net9764 net9896 vdd vss unit_coupling_tile
xi2395 net9893 net9693 net9904 net9894 net9891 net9901 net9692 net9892 vdd vss unit_coupling_tile
xi2394 net9903 net9689 net9905 net9904 net9901 net9899 net9688 net9902 vdd vss unit_coupling_tile
xi2393 net9912 net9699 net9909 net9905 net9899 net9906 net9698 net9900 vdd vss unit_coupling_tile
xi2392 net9908 net9708 net9910 net9909 net9906 net9911 net9696 net9907 vdd vss unit_coupling_tile
xi2391 net9917 net9704 net9918 net9910 net9911 net9913 net9703 net9916 vdd vss unit_coupling_tile
xi2390 net9915 net9713 net9922 net9918 net9913 net9919 net9712 net9914 vdd vss unit_coupling_tile
xi2389 net9921 net9711 net9923 net9922 net9919 net9924 net9710 net9920 vdd vss unit_coupling_tile
xi2388 net9930 net9717 net9928 net9923 net9924 net9925 net9716 net9929 vdd vss unit_coupling_tile
xi2387 net9927 net9726 net9857 net9928 net9925 net9931 net9725 net9926 vdd vss unit_coupling_tile
xi2386 net9856 net9723 net9853 net9857 net9931 net9850 net9722 net9932 vdd vss unit_coupling_tile
xi2385 net9852 net9652 net9854 net9853 net9850 net9855 net9728 net9851 vdd vss unit_coupling_tile
xi2384 net9862 net9648 net9863 net9854 net9855 net9858 net9647 net9861 vdd vss unit_coupling_tile
xi2383 net9860 net9658 net9867 net9863 net9858 net9864 net9657 net9859 vdd vss unit_coupling_tile
xi2382 net9866 net9656 net9868 net9867 net9864 net9869 net9655 net9865 vdd vss unit_coupling_tile
xi2381 net9875 net9662 net9873 net9868 net9869 net9870 net9661 net9874 vdd vss unit_coupling_tile
xi2380 net9872 net9671 net9881 net9873 net9870 net9878 net9670 net9871 vdd vss unit_coupling_tile
xi2379 net9880 net9668 net9882 net9881 net9878 net9876 net9667 net9879 vdd vss unit_coupling_tile
xi2378 net9888 net9676 net9886 net9882 net9876 net9883 net9675 net9877 vdd vss unit_coupling_tile
xi2377 net9885 net9684 net9815 net9886 net9883 net9887 net9673 net9884 vdd vss unit_coupling_tile
xi2376 net9890 net9681 net9812 net9815 net9887 net9809 net9680 net9889 vdd vss unit_coupling_tile
xi2375 net9811 net9686 net9813 net9812 net9809 net9814 net9685 net9810 vdd vss unit_coupling_tile
xi2374 net9821 net9607 net9819 net9813 net9814 net9816 net9606 net9820 vdd vss unit_coupling_tile
xi2373 net9818 net9617 net9827 net9819 net9816 net9824 net9616 net9817 vdd vss unit_coupling_tile
xi2372 net9826 net9614 net9828 net9827 net9824 net9822 net9613 net9825 vdd vss unit_coupling_tile
xi2371 net9835 net9622 net9832 net9828 net9822 net9829 net9621 net9823 vdd vss unit_coupling_tile
xi2370 net9831 net9631 net9833 net9832 net9829 net9834 net9619 net9830 vdd vss unit_coupling_tile
xi2369 net9840 net9627 net9841 net9833 net9834 net9836 net9626 net9839 vdd vss unit_coupling_tile
xi2368 net9838 net9636 net9845 net9841 net9836 net9842 net9635 net9837 vdd vss unit_coupling_tile
xi2367 net9844 net9634 net9846 net9845 net9842 net9847 net9633 net9843 vdd vss unit_coupling_tile
xi2366 net9849 net9640 net9774 net9846 net9847 net9771 net9639 net9848 vdd vss unit_coupling_tile
xi2365 net9773 net9645 net9775 net9774 net9771 net9769 net9644 net9772 vdd vss unit_coupling_tile
xi2364 net9782 net9569 net9779 net9775 net9769 net9776 net9568 net9770 vdd vss unit_coupling_tile
xi2363 net9778 net9578 net9780 net9779 net9776 net9781 net9566 net9777 vdd vss unit_coupling_tile
xi2362 net9787 net9574 net9788 net9780 net9781 net9783 net9573 net9786 vdd vss unit_coupling_tile
xi2361 net9785 net9583 net9792 net9788 net9783 net9789 net9582 net9784 vdd vss unit_coupling_tile
xi2360 net9791 net9581 net9793 net9792 net9789 net9794 net9580 net9790 vdd vss unit_coupling_tile
xi2359 net9800 net9587 net9798 net9793 net9794 net9795 net9586 net9799 vdd vss unit_coupling_tile
xi2358 net9797 net9596 net9806 net9798 net9795 net9803 net9595 net9796 vdd vss unit_coupling_tile
xi2357 net9805 net9593 net9807 net9806 net9803 net9801 net9592 net9804 vdd vss unit_coupling_tile
xi2356 net9808 net9601 net9735 net9807 net9801 net9732 net9600 net9802 vdd vss unit_coupling_tile
xi2355 net9734 net9604 net9736 net9735 net9732 net9729 net9598 net9733 vdd vss unit_coupling_tile
xi2354 net9731 net9527 net9740 net9736 net9729 net9737 net9526 net9730 vdd vss unit_coupling_tile
xi2353 net9739 net9532 net9741 net9740 net9737 net9742 net9531 net9738 vdd vss unit_coupling_tile
xi2351 net9745 net9544 net9753 net9746 net9743 net9750 net9543 net9744 vdd vss unit_coupling_tile
xi2350 net9752 net9541 net9754 net9753 net9750 net9755 net9540 net9751 vdd vss unit_coupling_tile
xi2349 net9762 net9548 net9759 net56 net56 net9756 net9547 net9749 vdd vss unit_coupling_tile
xi2348 net9758 net9558 net9760 net9759 net9756 net9761 net9546 net9757 vdd vss unit_coupling_tile
xi2347 net9767 net9554 net9768 net9760 net9761 net9763 net9553 net9766 vdd vss unit_coupling_tile
xi2346 net9765 net9563 net9694 net9768 net9763 net9691 net9562 net9764 vdd vss unit_coupling_tile
xi2345 net9693 net9561 net9690 net9694 net9691 net9687 net9560 net9692 vdd vss unit_coupling_tile
xi2344 net9689 net9489 net9700 net9690 net9687 net9697 net9488 net9688 vdd vss unit_coupling_tile
xi2343 net9699 net9485 net9701 net9700 net9697 net9695 net9484 net9698 vdd vss unit_coupling_tile
xi2342 net9708 net9495 net9705 net9701 net9695 net9702 net9494 net9696 vdd vss unit_coupling_tile
xi2341 net9704 net9504 net9706 net9705 net9702 net9707 net9492 net9703 vdd vss unit_coupling_tile
xi2340 net9713 net9500 net9714 net9706 net9707 net9709 net9499 net9712 vdd vss unit_coupling_tile
xi2339 net9711 net9509 net9718 net9714 net9709 net9715 net9508 net9710 vdd vss unit_coupling_tile
xi2338 net9717 net9507 net9719 net9718 net9715 net9720 net9506 net9716 vdd vss unit_coupling_tile
xi2337 net9726 net9513 net9724 net9719 net9720 net9721 net9512 net9725 vdd vss unit_coupling_tile
xi2336 net9723 net9522 net9653 net9724 net9721 net9727 net9521 net9722 vdd vss unit_coupling_tile
xi2335 net9652 net9519 net9649 net9653 net9727 net9646 net9518 net9728 vdd vss unit_coupling_tile
xi2334 net9648 net9448 net9650 net9649 net9646 net9651 net9524 net9647 vdd vss unit_coupling_tile
xi2333 net9658 net9444 net9659 net9650 net9651 net9654 net9443 net9657 vdd vss unit_coupling_tile
xi2332 net9656 net9454 net9663 net9659 net9654 net9660 net9453 net9655 vdd vss unit_coupling_tile
xi2331 net9662 net9452 net9664 net9663 net9660 net9665 net9451 net9661 vdd vss unit_coupling_tile
xi2330 net9671 net9458 net9669 net9664 net9665 net9666 net9457 net9670 vdd vss unit_coupling_tile
xi2329 net9668 net9467 net9677 net9669 net9666 net9674 net9466 net9667 vdd vss unit_coupling_tile
xi2328 net9676 net9464 net9678 net9677 net9674 net9672 net9463 net9675 vdd vss unit_coupling_tile
xi2327 net9684 net9472 net9682 net9678 net9672 net9679 net9471 net9673 vdd vss unit_coupling_tile
xi2326 net9681 net9480 net9611 net9682 net9679 net9683 net9469 net9680 vdd vss unit_coupling_tile
xi2325 net9686 net9477 net9608 net9611 net9683 net9605 net9476 net9685 vdd vss unit_coupling_tile
xi2324 net9607 net9482 net9609 net9608 net9605 net9610 net9481 net9606 vdd vss unit_coupling_tile
xi2323 net9617 net9403 net9615 net9609 net9610 net9612 net9402 net9616 vdd vss unit_coupling_tile
xi2322 net9614 net9413 net9623 net9615 net9612 net9620 net9412 net9613 vdd vss unit_coupling_tile
xi2321 net9622 net9410 net9624 net9623 net9620 net9618 net9409 net9621 vdd vss unit_coupling_tile
xi2320 net9631 net9418 net9628 net9624 net9618 net9625 net9417 net9619 vdd vss unit_coupling_tile
xi2319 net9627 net9427 net9629 net9628 net9625 net9630 net9415 net9626 vdd vss unit_coupling_tile
xi2318 net9636 net9423 net9637 net9629 net9630 net9632 net9422 net9635 vdd vss unit_coupling_tile
xi2317 net9634 net9432 net9641 net9637 net9632 net9638 net9431 net9633 vdd vss unit_coupling_tile
xi2316 net9640 net9430 net9642 net9641 net9638 net9643 net9429 net9639 vdd vss unit_coupling_tile
xi2315 net9645 net9436 net9570 net9642 net9643 net9567 net9435 net9644 vdd vss unit_coupling_tile
xi2314 net9569 net9441 net9571 net9570 net9567 net9565 net9440 net9568 vdd vss unit_coupling_tile
xi2313 net9578 net9365 net9575 net9571 net9565 net9572 net9364 net9566 vdd vss unit_coupling_tile
xi2312 net9574 net9374 net9576 net9575 net9572 net9577 net9362 net9573 vdd vss unit_coupling_tile
xi2311 net9583 net9370 net9584 net9576 net9577 net9579 net9369 net9582 vdd vss unit_coupling_tile
xi2310 net9581 net9379 net9588 net9584 net9579 net9585 net9378 net9580 vdd vss unit_coupling_tile
xi2309 net9587 net9377 net9589 net9588 net9585 net9590 net9376 net9586 vdd vss unit_coupling_tile
xi2308 net9596 net9383 net9594 net9589 net9590 net9591 net9382 net9595 vdd vss unit_coupling_tile
xi2307 net9593 net9392 net9602 net9594 net9591 net9599 net9391 net9592 vdd vss unit_coupling_tile
xi2306 net9601 net9389 net9603 net9602 net9599 net9597 net9388 net9600 vdd vss unit_coupling_tile
xi2305 net9604 net9395 net9528 net9603 net9597 net9525 net9394 net9598 vdd vss unit_coupling_tile
xi2304 net9527 net9400 net9529 net9528 net9525 net9530 net9399 net9526 vdd vss unit_coupling_tile
xi2302 net9535 net9323 net9537 net9536 net9533 net9538 net9322 net9534 vdd vss unit_coupling_tile
xi2301 net9544 net9331 net9542 net9537 net9538 net9539 net9330 net9543 vdd vss unit_coupling_tile
xi2300 net9541 net9338 net9550 net9542 net9539 net9551 net9337 net9540 vdd vss unit_coupling_tile
xi2299 net9548 net9336 net9549 net57 net57 net9545 net9335 net9547 vdd vss unit_coupling_tile
xi2298 net9558 net9345 net9555 net9549 net9545 net9552 net9344 net9546 vdd vss unit_coupling_tile
xi2297 net9554 net9354 net9556 net9555 net9552 net9557 net9342 net9553 vdd vss unit_coupling_tile
xi2296 net9563 net9350 net9564 net9556 net9557 net9559 net9349 net9562 vdd vss unit_coupling_tile
xi2295 net9561 net9359 net9490 net9564 net9559 net9487 net9358 net9560 vdd vss unit_coupling_tile
xi2294 net9489 net9357 net9486 net9490 net9487 net9483 net9356 net9488 vdd vss unit_coupling_tile
xi2293 net9485 net9285 net9496 net9486 net9483 net9493 net9284 net9484 vdd vss unit_coupling_tile
xi2292 net9495 net9281 net9497 net9496 net9493 net9491 net9280 net9494 vdd vss unit_coupling_tile
xi2291 net9504 net9291 net9501 net9497 net9491 net9498 net9290 net9492 vdd vss unit_coupling_tile
xi2290 net9500 net9300 net9502 net9501 net9498 net9503 net9288 net9499 vdd vss unit_coupling_tile
xi2289 net9509 net9296 net9510 net9502 net9503 net9505 net9295 net9508 vdd vss unit_coupling_tile
xi2288 net9507 net9305 net9514 net9510 net9505 net9511 net9304 net9506 vdd vss unit_coupling_tile
xi2287 net9513 net9303 net9515 net9514 net9511 net9516 net9302 net9512 vdd vss unit_coupling_tile
xi2286 net9522 net9309 net9520 net9515 net9516 net9517 net9308 net9521 vdd vss unit_coupling_tile
xi2285 net9519 net9318 net9449 net9520 net9517 net9523 net9317 net9518 vdd vss unit_coupling_tile
xi2284 net9448 net9315 net9445 net9449 net9523 net9442 net9314 net9524 vdd vss unit_coupling_tile
xi2283 net9444 net9244 net9446 net9445 net9442 net9447 net9320 net9443 vdd vss unit_coupling_tile
xi2282 net9454 net9240 net9455 net9446 net9447 net9450 net9239 net9453 vdd vss unit_coupling_tile
xi2281 net9452 net9250 net9459 net9455 net9450 net9456 net9249 net9451 vdd vss unit_coupling_tile
xi2280 net9458 net9248 net9460 net9459 net9456 net9461 net9247 net9457 vdd vss unit_coupling_tile
xi2279 net9467 net9254 net9465 net9460 net9461 net9462 net9253 net9466 vdd vss unit_coupling_tile
xi2278 net9464 net9263 net9473 net9465 net9462 net9470 net9262 net9463 vdd vss unit_coupling_tile
xi2277 net9472 net9260 net9474 net9473 net9470 net9468 net9259 net9471 vdd vss unit_coupling_tile
xi2276 net9480 net9268 net9478 net9474 net9468 net9475 net9267 net9469 vdd vss unit_coupling_tile
xi2275 net9477 net9276 net9407 net9478 net9475 net9479 net9265 net9476 vdd vss unit_coupling_tile
xi2274 net9482 net9273 net9404 net9407 net9479 net9401 net9272 net9481 vdd vss unit_coupling_tile
xi2273 net9403 net9278 net9405 net9404 net9401 net9406 net9277 net9402 vdd vss unit_coupling_tile
xi2272 net9413 net9199 net9411 net9405 net9406 net9408 net9198 net9412 vdd vss unit_coupling_tile
xi2271 net9410 net9209 net9419 net9411 net9408 net9416 net9208 net9409 vdd vss unit_coupling_tile
xi2270 net9418 net9206 net9420 net9419 net9416 net9414 net9205 net9417 vdd vss unit_coupling_tile
xi2269 net9427 net9214 net9424 net9420 net9414 net9421 net9213 net9415 vdd vss unit_coupling_tile
xi2268 net9423 net9223 net9425 net9424 net9421 net9426 net9211 net9422 vdd vss unit_coupling_tile
xi2267 net9432 net9219 net9433 net9425 net9426 net9428 net9218 net9431 vdd vss unit_coupling_tile
xi2266 net9430 net9228 net9437 net9433 net9428 net9434 net9227 net9429 vdd vss unit_coupling_tile
xi2265 net9436 net9226 net9438 net9437 net9434 net9439 net9225 net9435 vdd vss unit_coupling_tile
xi2264 net9441 net9232 net9366 net9438 net9439 net9363 net9231 net9440 vdd vss unit_coupling_tile
xi2263 net9365 net9237 net9367 net9366 net9363 net9361 net9236 net9364 vdd vss unit_coupling_tile
xi2262 net9374 net9161 net9371 net9367 net9361 net9368 net9160 net9362 vdd vss unit_coupling_tile
xi2261 net9370 net9170 net9372 net9371 net9368 net9373 net9158 net9369 vdd vss unit_coupling_tile
xi2260 net9379 net9166 net9380 net9372 net9373 net9375 net9165 net9378 vdd vss unit_coupling_tile
xi2259 net9377 net9175 net9384 net9380 net9375 net9381 net9174 net9376 vdd vss unit_coupling_tile
xi2258 net9383 net9173 net9385 net9384 net9381 net9386 net9172 net9382 vdd vss unit_coupling_tile
xi2257 net9392 net9179 net9390 net9385 net9386 net9387 net9178 net9391 vdd vss unit_coupling_tile
xi2256 net9389 net9184 net9396 net9390 net9387 net9393 net9183 net9388 vdd vss unit_coupling_tile
xi2255 net9395 net9188 net9397 net9396 net9393 net9398 net9187 net9394 vdd vss unit_coupling_tile
xi2253 net9326 net9196 net9328 net9327 net9324 net9321 net9190 net9325 vdd vss unit_coupling_tile
xi2252 net9323 net9122 net9332 net9328 net9321 net9329 net9121 net9322 vdd vss unit_coupling_tile
xi2251 net9331 net9119 net9333 net9332 net9329 net9334 net9118 net9330 vdd vss unit_coupling_tile
xi2250 net9338 net9127 net9339 net9333 net9334 net9340 net9126 net9337 vdd vss unit_coupling_tile
xi2249 net9336 net9136 net9346 net58 net58 net9343 net9135 net9335 vdd vss unit_coupling_tile
xi2248 net9345 net9133 net9347 net9346 net9343 net9341 net9132 net9344 vdd vss unit_coupling_tile
xi2247 net9354 net9141 net9351 net9347 net9341 net9348 net9140 net9342 vdd vss unit_coupling_tile
xi2246 net9350 net9150 net9352 net9351 net9348 net9353 net9138 net9349 vdd vss unit_coupling_tile
xi2245 net9359 net9146 net9360 net9352 net9353 net9355 net9145 net9358 vdd vss unit_coupling_tile
xi2244 net9357 net9155 net9286 net9360 net9355 net9283 net9154 net9356 vdd vss unit_coupling_tile
xi2243 net9285 net9153 net9282 net9286 net9283 net9279 net9152 net9284 vdd vss unit_coupling_tile
xi2242 net9281 net9081 net9292 net9282 net9279 net9289 net9080 net9280 vdd vss unit_coupling_tile
xi2241 net9291 net9077 net9293 net9292 net9289 net9287 net9076 net9290 vdd vss unit_coupling_tile
xi2240 net9300 net9087 net9297 net9293 net9287 net9294 net9086 net9288 vdd vss unit_coupling_tile
xi2239 net9296 net9096 net9298 net9297 net9294 net9299 net9084 net9295 vdd vss unit_coupling_tile
xi2238 net9305 net9092 net9306 net9298 net9299 net9301 net9091 net9304 vdd vss unit_coupling_tile
xi2237 net9303 net9101 net9310 net9306 net9301 net9307 net9100 net9302 vdd vss unit_coupling_tile
xi2236 net9309 net9099 net9311 net9310 net9307 net9312 net9098 net9308 vdd vss unit_coupling_tile
xi2235 net9318 net9105 net9316 net9311 net9312 net9313 net9104 net9317 vdd vss unit_coupling_tile
xi2234 net9315 net9114 net9245 net9316 net9313 net9319 net9113 net9314 vdd vss unit_coupling_tile
xi2233 net9244 net9111 net9241 net9245 net9319 net9238 net9110 net9320 vdd vss unit_coupling_tile
xi2232 net9240 net9040 net9242 net9241 net9238 net9243 net9116 net9239 vdd vss unit_coupling_tile
xi2231 net9250 net9036 net9251 net9242 net9243 net9246 net9035 net9249 vdd vss unit_coupling_tile
xi2230 net9248 net9046 net9255 net9251 net9246 net9252 net9045 net9247 vdd vss unit_coupling_tile
xi2229 net9254 net9044 net9256 net9255 net9252 net9257 net9043 net9253 vdd vss unit_coupling_tile
xi2228 net9263 net9050 net9261 net9256 net9257 net9258 net9049 net9262 vdd vss unit_coupling_tile
xi2227 net9260 net9059 net9269 net9261 net9258 net9266 net9058 net9259 vdd vss unit_coupling_tile
xi2226 net9268 net9056 net9270 net9269 net9266 net9264 net9055 net9267 vdd vss unit_coupling_tile
xi2225 net9276 net9064 net9274 net9270 net9264 net9271 net9063 net9265 vdd vss unit_coupling_tile
xi2224 net9273 net9072 net9203 net9274 net9271 net9275 net9061 net9272 vdd vss unit_coupling_tile
xi2223 net9278 net9069 net9200 net9203 net9275 net9197 net9068 net9277 vdd vss unit_coupling_tile
xi2222 net9199 net9074 net9201 net9200 net9197 net9202 net9073 net9198 vdd vss unit_coupling_tile
xi2221 net9209 net8995 net9207 net9201 net9202 net9204 net8994 net9208 vdd vss unit_coupling_tile
xi2220 net9206 net9005 net9215 net9207 net9204 net9212 net9004 net9205 vdd vss unit_coupling_tile
xi2219 net9214 net9002 net9216 net9215 net9212 net9210 net9001 net9213 vdd vss unit_coupling_tile
xi2218 net9223 net9010 net9220 net9216 net9210 net9217 net9009 net9211 vdd vss unit_coupling_tile
xi2217 net9219 net9019 net9221 net9220 net9217 net9222 net9007 net9218 vdd vss unit_coupling_tile
xi2216 net9228 net9015 net9229 net9221 net9222 net9224 net9014 net9227 vdd vss unit_coupling_tile
xi2215 net9226 net9024 net9233 net9229 net9224 net9230 net9023 net9225 vdd vss unit_coupling_tile
xi2214 net9232 net9022 net9234 net9233 net9230 net9235 net9021 net9231 vdd vss unit_coupling_tile
xi2213 net9237 net9028 net9162 net9234 net9235 net9159 net9027 net9236 vdd vss unit_coupling_tile
xi2212 net9161 net9033 net9163 net9162 net9159 net9157 net9032 net9160 vdd vss unit_coupling_tile
xi2211 net9170 net8957 net9167 net9163 net9157 net9164 net8956 net9158 vdd vss unit_coupling_tile
xi2210 net9166 net8966 net9168 net9167 net9164 net9169 net8954 net9165 vdd vss unit_coupling_tile
xi2209 net9175 net8962 net9176 net9168 net9169 net9171 net8961 net9174 vdd vss unit_coupling_tile
xi2208 net9173 net8971 net9180 net9176 net9171 net9177 net8970 net9172 vdd vss unit_coupling_tile
xi2207 net9179 net8969 net9181 net9180 net9177 net9182 net8968 net9178 vdd vss unit_coupling_tile
xi2206 net9184 net8976 net9185 net9181 net9182 net9186 net8975 net9183 vdd vss unit_coupling_tile
xi2204 net9193 net8981 net9195 net9194 net9191 net9189 net8980 net9192 vdd vss unit_coupling_tile
xi2203 net9196 net8989 net9123 net9195 net9189 net9120 net8988 net9190 vdd vss unit_coupling_tile
xi2202 net9122 net8992 net9124 net9123 net9120 net9117 net8986 net9121 vdd vss unit_coupling_tile
xi2201 net9119 net8918 net9128 net9124 net9117 net9125 net8917 net9118 vdd vss unit_coupling_tile
xi2200 net9127 net8915 net9129 net9128 net9125 net9130 net8914 net9126 vdd vss unit_coupling_tile
xi2199 net9136 net8922 net9134 net59 net59 net9131 net8921 net9135 vdd vss unit_coupling_tile
xi2198 net9133 net8932 net9142 net9134 net9131 net9139 net8931 net9132 vdd vss unit_coupling_tile
xi2197 net9141 net8929 net9143 net9142 net9139 net9137 net8928 net9140 vdd vss unit_coupling_tile
xi2196 net9150 net8937 net9147 net9143 net9137 net9144 net8936 net9138 vdd vss unit_coupling_tile
xi2195 net9146 net8946 net9148 net9147 net9144 net9149 net8934 net9145 vdd vss unit_coupling_tile
xi2194 net9155 net8942 net9156 net9148 net9149 net9151 net8941 net9154 vdd vss unit_coupling_tile
xi2193 net9153 net8951 net9082 net9156 net9151 net9079 net8950 net9152 vdd vss unit_coupling_tile
xi2192 net9081 net8949 net9078 net9082 net9079 net9075 net8948 net9080 vdd vss unit_coupling_tile
xi2191 net9077 net8877 net9088 net9078 net9075 net9085 net8876 net9076 vdd vss unit_coupling_tile
xi2190 net9087 net8873 net9089 net9088 net9085 net9083 net8872 net9086 vdd vss unit_coupling_tile
xi2189 net9096 net8883 net9093 net9089 net9083 net9090 net8882 net9084 vdd vss unit_coupling_tile
xi2188 net9092 net8892 net9094 net9093 net9090 net9095 net8880 net9091 vdd vss unit_coupling_tile
xi2187 net9101 net8888 net9102 net9094 net9095 net9097 net8887 net9100 vdd vss unit_coupling_tile
xi2186 net9099 net8897 net9106 net9102 net9097 net9103 net8896 net9098 vdd vss unit_coupling_tile
xi2185 net9105 net8895 net9107 net9106 net9103 net9108 net8894 net9104 vdd vss unit_coupling_tile
xi2184 net9114 net8901 net9112 net9107 net9108 net9109 net8900 net9113 vdd vss unit_coupling_tile
xi2183 net9111 net8910 net9041 net9112 net9109 net9115 net8909 net9110 vdd vss unit_coupling_tile
xi2182 net9040 net8907 net9037 net9041 net9115 net9034 net8906 net9116 vdd vss unit_coupling_tile
xi2181 net9036 net8836 net9038 net9037 net9034 net9039 net8912 net9035 vdd vss unit_coupling_tile
xi2180 net9046 net8832 net9047 net9038 net9039 net9042 net8831 net9045 vdd vss unit_coupling_tile
xi2179 net9044 net8842 net9051 net9047 net9042 net9048 net8841 net9043 vdd vss unit_coupling_tile
xi2178 net9050 net8840 net9052 net9051 net9048 net9053 net8839 net9049 vdd vss unit_coupling_tile
xi2177 net9059 net8846 net9057 net9052 net9053 net9054 net8845 net9058 vdd vss unit_coupling_tile
xi2176 net9056 net8855 net9065 net9057 net9054 net9062 net8854 net9055 vdd vss unit_coupling_tile
xi2175 net9064 net8852 net9066 net9065 net9062 net9060 net8851 net9063 vdd vss unit_coupling_tile
xi2174 net9072 net8860 net9070 net9066 net9060 net9067 net8859 net9061 vdd vss unit_coupling_tile
xi2173 net9069 net8868 net8999 net9070 net9067 net9071 net8857 net9068 vdd vss unit_coupling_tile
xi2172 net9074 net8865 net8996 net8999 net9071 net8993 net8864 net9073 vdd vss unit_coupling_tile
xi2171 net8995 net8870 net8997 net8996 net8993 net8998 net8869 net8994 vdd vss unit_coupling_tile
xi2170 net9005 net8791 net9003 net8997 net8998 net9000 net8790 net9004 vdd vss unit_coupling_tile
xi2169 net9002 net8801 net9011 net9003 net9000 net9008 net8800 net9001 vdd vss unit_coupling_tile
xi2168 net9010 net8798 net9012 net9011 net9008 net9006 net8797 net9009 vdd vss unit_coupling_tile
xi2167 net9019 net8806 net9016 net9012 net9006 net9013 net8805 net9007 vdd vss unit_coupling_tile
xi2166 net9015 net8815 net9017 net9016 net9013 net9018 net8803 net9014 vdd vss unit_coupling_tile
xi2165 net9024 net8811 net9025 net9017 net9018 net9020 net8810 net9023 vdd vss unit_coupling_tile
xi2164 net9022 net8820 net9029 net9025 net9020 net9026 net8819 net9021 vdd vss unit_coupling_tile
xi2163 net9028 net8818 net9030 net9029 net9026 net9031 net8817 net9027 vdd vss unit_coupling_tile
xi2162 net9033 net8824 net8958 net9030 net9031 net8955 net8823 net9032 vdd vss unit_coupling_tile
xi2161 net8957 net8829 net8959 net8958 net8955 net8953 net8828 net8956 vdd vss unit_coupling_tile
xi2160 net8966 net8753 net8963 net8959 net8953 net8960 net8752 net8954 vdd vss unit_coupling_tile
xi2159 net8962 net8762 net8964 net8963 net8960 net8965 net8750 net8961 vdd vss unit_coupling_tile
xi2158 net8971 net8758 net8972 net8964 net8965 net8967 net8757 net8970 vdd vss unit_coupling_tile
xi2157 net8969 net8767 net8973 net8972 net8967 net8974 net8766 net8968 vdd vss unit_coupling_tile
xi2155 net8984 net8771 net8982 net8977 net8978 net8979 net8770 net8983 vdd vss unit_coupling_tile
xi2154 net8981 net8780 net8990 net8982 net8979 net8987 net8779 net8980 vdd vss unit_coupling_tile
xi2153 net8989 net8777 net8991 net8990 net8987 net8985 net8776 net8988 vdd vss unit_coupling_tile
xi2152 net8992 net8785 net8919 net8991 net8985 net8916 net8784 net8986 vdd vss unit_coupling_tile
xi2151 net8918 net8788 net8920 net8919 net8916 net8913 net8782 net8917 vdd vss unit_coupling_tile
xi2150 net8915 net8713 net8925 net8920 net8913 net8926 net8712 net8914 vdd vss unit_coupling_tile
xi2149 net8922 net8710 net8923 net60 net60 net8924 net8709 net8921 vdd vss unit_coupling_tile
xi2148 net8932 net8719 net8930 net8923 net8924 net8927 net8718 net8931 vdd vss unit_coupling_tile
xi2147 net8929 net8728 net8938 net8930 net8927 net8935 net8727 net8928 vdd vss unit_coupling_tile
xi2146 net8937 net8725 net8939 net8938 net8935 net8933 net8724 net8936 vdd vss unit_coupling_tile
xi2145 net8946 net8733 net8943 net8939 net8933 net8940 net8732 net8934 vdd vss unit_coupling_tile
xi2144 net8942 net8742 net8944 net8943 net8940 net8945 net8730 net8941 vdd vss unit_coupling_tile
xi2143 net8951 net8738 net8952 net8944 net8945 net8947 net8737 net8950 vdd vss unit_coupling_tile
xi2142 net8949 net8747 net8878 net8952 net8947 net8875 net8746 net8948 vdd vss unit_coupling_tile
xi2141 net8877 net8745 net8874 net8878 net8875 net8871 net8744 net8876 vdd vss unit_coupling_tile
xi2140 net8873 net8673 net8884 net8874 net8871 net8881 net8672 net8872 vdd vss unit_coupling_tile
xi2139 net8883 net8669 net8885 net8884 net8881 net8879 net8668 net8882 vdd vss unit_coupling_tile
xi2138 net8892 net8679 net8889 net8885 net8879 net8886 net8678 net8880 vdd vss unit_coupling_tile
xi2137 net8888 net8688 net8890 net8889 net8886 net8891 net8676 net8887 vdd vss unit_coupling_tile
xi2136 net8897 net8684 net8898 net8890 net8891 net8893 net8683 net8896 vdd vss unit_coupling_tile
xi2135 net8895 net8693 net8902 net8898 net8893 net8899 net8692 net8894 vdd vss unit_coupling_tile
xi2134 net8901 net8691 net8903 net8902 net8899 net8904 net8690 net8900 vdd vss unit_coupling_tile
xi2133 net8910 net8697 net8908 net8903 net8904 net8905 net8696 net8909 vdd vss unit_coupling_tile
xi2132 net8907 net8706 net8837 net8908 net8905 net8911 net8705 net8906 vdd vss unit_coupling_tile
xi2131 net8836 net8703 net8833 net8837 net8911 net8830 net8702 net8912 vdd vss unit_coupling_tile
xi2130 net8832 net8632 net8834 net8833 net8830 net8835 net8708 net8831 vdd vss unit_coupling_tile
xi2129 net8842 net8628 net8843 net8834 net8835 net8838 net8627 net8841 vdd vss unit_coupling_tile
xi2128 net8840 net8638 net8847 net8843 net8838 net8844 net8637 net8839 vdd vss unit_coupling_tile
xi2127 net8846 net8636 net8848 net8847 net8844 net8849 net8635 net8845 vdd vss unit_coupling_tile
xi2126 net8855 net8642 net8853 net8848 net8849 net8850 net8641 net8854 vdd vss unit_coupling_tile
xi2125 net8852 net8651 net8861 net8853 net8850 net8858 net8650 net8851 vdd vss unit_coupling_tile
xi2124 net8860 net8648 net8862 net8861 net8858 net8856 net8647 net8859 vdd vss unit_coupling_tile
xi2123 net8868 net8656 net8866 net8862 net8856 net8863 net8655 net8857 vdd vss unit_coupling_tile
xi2122 net8865 net8664 net8795 net8866 net8863 net8867 net8653 net8864 vdd vss unit_coupling_tile
xi2121 net8870 net8661 net8792 net8795 net8867 net8789 net8660 net8869 vdd vss unit_coupling_tile
xi2120 net8791 net8666 net8793 net8792 net8789 net8794 net8665 net8790 vdd vss unit_coupling_tile
xi2119 net8801 net8587 net8799 net8793 net8794 net8796 net8586 net8800 vdd vss unit_coupling_tile
xi2118 net8798 net8597 net8807 net8799 net8796 net8804 net8596 net8797 vdd vss unit_coupling_tile
xi2117 net8806 net8594 net8808 net8807 net8804 net8802 net8593 net8805 vdd vss unit_coupling_tile
xi2116 net8815 net8602 net8812 net8808 net8802 net8809 net8601 net8803 vdd vss unit_coupling_tile
xi2115 net8811 net8611 net8813 net8812 net8809 net8814 net8599 net8810 vdd vss unit_coupling_tile
xi2114 net8820 net8607 net8821 net8813 net8814 net8816 net8606 net8819 vdd vss unit_coupling_tile
xi2113 net8818 net8616 net8825 net8821 net8816 net8822 net8615 net8817 vdd vss unit_coupling_tile
xi2112 net8824 net8614 net8826 net8825 net8822 net8827 net8613 net8823 vdd vss unit_coupling_tile
xi2111 net8829 net8620 net8754 net8826 net8827 net8751 net8619 net8828 vdd vss unit_coupling_tile
xi2110 net8753 net8625 net8755 net8754 net8751 net8749 net8624 net8752 vdd vss unit_coupling_tile
xi2109 net8762 net8545 net8759 net8755 net8749 net8756 net8544 net8750 vdd vss unit_coupling_tile
xi2108 net8758 net8556 net8760 net8759 net8756 net8761 net8549 net8757 vdd vss unit_coupling_tile
xi2106 net8765 net8561 net8772 net8768 net8763 net8769 net8560 net8764 vdd vss unit_coupling_tile
xi2105 net8771 net8559 net8773 net8772 net8769 net8774 net8558 net8770 vdd vss unit_coupling_tile
xi2104 net8780 net8565 net8778 net8773 net8774 net8775 net8564 net8779 vdd vss unit_coupling_tile
xi2103 net8777 net8574 net8786 net8778 net8775 net8783 net8573 net8776 vdd vss unit_coupling_tile
xi2102 net8785 net8571 net8787 net8786 net8783 net8781 net8570 net8784 vdd vss unit_coupling_tile
xi2101 net8788 net8579 net8714 net8787 net8781 net8711 net8578 net8782 vdd vss unit_coupling_tile
xi2100 net8713 net8582 net8715 net8714 net8711 net8716 net8576 net8712 vdd vss unit_coupling_tile
xi2099 net8710 net8509 net8720 net61 net61 net8717 net8508 net8709 vdd vss unit_coupling_tile
xi2098 net8719 net8507 net8721 net8720 net8717 net8722 net8506 net8718 vdd vss unit_coupling_tile
xi2097 net8728 net8513 net8726 net8721 net8722 net8723 net8512 net8727 vdd vss unit_coupling_tile
xi2096 net8725 net8522 net8734 net8726 net8723 net8731 net8521 net8724 vdd vss unit_coupling_tile
xi2095 net8733 net8519 net8735 net8734 net8731 net8729 net8518 net8732 vdd vss unit_coupling_tile
xi2094 net8742 net8527 net8739 net8735 net8729 net8736 net8526 net8730 vdd vss unit_coupling_tile
xi2093 net8738 net8536 net8740 net8739 net8736 net8741 net8524 net8737 vdd vss unit_coupling_tile
xi2092 net8747 net8532 net8748 net8740 net8741 net8743 net8531 net8746 vdd vss unit_coupling_tile
xi2091 net8745 net8541 net8674 net8748 net8743 net8671 net8540 net8744 vdd vss unit_coupling_tile
xi2090 net8673 net8539 net8670 net8674 net8671 net8667 net8538 net8672 vdd vss unit_coupling_tile
xi2089 net8669 net8469 net8680 net8670 net8667 net8677 net8468 net8668 vdd vss unit_coupling_tile
xi2088 net8679 net8465 net8681 net8680 net8677 net8675 net8464 net8678 vdd vss unit_coupling_tile
xi2087 net8688 net8475 net8685 net8681 net8675 net8682 net8474 net8676 vdd vss unit_coupling_tile
xi2086 net8684 net8484 net8686 net8685 net8682 net8687 net8472 net8683 vdd vss unit_coupling_tile
xi2085 net8693 net8480 net8694 net8686 net8687 net8689 net8479 net8692 vdd vss unit_coupling_tile
xi2084 net8691 net8489 net8698 net8694 net8689 net8695 net8488 net8690 vdd vss unit_coupling_tile
xi2083 net8697 net8487 net8699 net8698 net8695 net8700 net8486 net8696 vdd vss unit_coupling_tile
xi2082 net8706 net8493 net8704 net8699 net8700 net8701 net8492 net8705 vdd vss unit_coupling_tile
xi2081 net8703 net8502 net8633 net8704 net8701 net8707 net8501 net8702 vdd vss unit_coupling_tile
xi2080 net8632 net8499 net8629 net8633 net8707 net8626 net8498 net8708 vdd vss unit_coupling_tile
xi2079 net8628 net8428 net8630 net8629 net8626 net8631 net8504 net8627 vdd vss unit_coupling_tile
xi2078 net8638 net8424 net8639 net8630 net8631 net8634 net8423 net8637 vdd vss unit_coupling_tile
xi2077 net8636 net8434 net8643 net8639 net8634 net8640 net8433 net8635 vdd vss unit_coupling_tile
xi2076 net8642 net8432 net8644 net8643 net8640 net8645 net8431 net8641 vdd vss unit_coupling_tile
xi2075 net8651 net8438 net8649 net8644 net8645 net8646 net8437 net8650 vdd vss unit_coupling_tile
xi2074 net8648 net8447 net8657 net8649 net8646 net8654 net8446 net8647 vdd vss unit_coupling_tile
xi2073 net8656 net8444 net8658 net8657 net8654 net8652 net8443 net8655 vdd vss unit_coupling_tile
xi2072 net8664 net8452 net8662 net8658 net8652 net8659 net8451 net8653 vdd vss unit_coupling_tile
xi2071 net8661 net8460 net8591 net8662 net8659 net8663 net8449 net8660 vdd vss unit_coupling_tile
xi2070 net8666 net8457 net8588 net8591 net8663 net8585 net8456 net8665 vdd vss unit_coupling_tile
xi2069 net8587 net8462 net8589 net8588 net8585 net8590 net8461 net8586 vdd vss unit_coupling_tile
xi2068 net8597 net8383 net8595 net8589 net8590 net8592 net8382 net8596 vdd vss unit_coupling_tile
xi2067 net8594 net8393 net8603 net8595 net8592 net8600 net8392 net8593 vdd vss unit_coupling_tile
xi2066 net8602 net8390 net8604 net8603 net8600 net8598 net8389 net8601 vdd vss unit_coupling_tile
xi2065 net8611 net8398 net8608 net8604 net8598 net8605 net8397 net8599 vdd vss unit_coupling_tile
xi2064 net8607 net8407 net8609 net8608 net8605 net8610 net8395 net8606 vdd vss unit_coupling_tile
xi2063 net8616 net8403 net8617 net8609 net8610 net8612 net8402 net8615 vdd vss unit_coupling_tile
xi2062 net8614 net8412 net8621 net8617 net8612 net8618 net8411 net8613 vdd vss unit_coupling_tile
xi2061 net8620 net8410 net8622 net8621 net8618 net8623 net8409 net8619 vdd vss unit_coupling_tile
xi2060 net8625 net8416 net8546 net8622 net8623 net8543 net8415 net8624 vdd vss unit_coupling_tile
xi2059 net8545 net8421 net8547 net8546 net8543 net8548 net8420 net8544 vdd vss unit_coupling_tile
xi2057 net8552 net8354 net8554 net8553 net8550 net8555 net8342 net8551 vdd vss unit_coupling_tile
xi2056 net8561 net8350 net8562 net8554 net8555 net8557 net8349 net8560 vdd vss unit_coupling_tile
xi2055 net8559 net8359 net8566 net8562 net8557 net8563 net8358 net8558 vdd vss unit_coupling_tile
xi2054 net8565 net8357 net8567 net8566 net8563 net8568 net8356 net8564 vdd vss unit_coupling_tile
xi2053 net8574 net8363 net8572 net8567 net8568 net8569 net8362 net8573 vdd vss unit_coupling_tile
xi2052 net8571 net8372 net8580 net8572 net8569 net8577 net8371 net8570 vdd vss unit_coupling_tile
xi2051 net8579 net8369 net8581 net8580 net8577 net8575 net8368 net8578 vdd vss unit_coupling_tile
xi2050 net8582 net8376 net8583 net8581 net8575 net8584 net8375 net8576 vdd vss unit_coupling_tile
xi2049 net8509 net8380 net8510 net62 net62 net8505 net8373 net8508 vdd vss unit_coupling_tile
xi2048 net8507 net8306 net8514 net8510 net8505 net8511 net8305 net8506 vdd vss unit_coupling_tile
xi2047 net8513 net8303 net8515 net8514 net8511 net8516 net8302 net8512 vdd vss unit_coupling_tile
xi2046 net8522 net8311 net8520 net8515 net8516 net8517 net8310 net8521 vdd vss unit_coupling_tile
xi2045 net8519 net8320 net8528 net8520 net8517 net8525 net8319 net8518 vdd vss unit_coupling_tile
xi2044 net8527 net8317 net8529 net8528 net8525 net8523 net8316 net8526 vdd vss unit_coupling_tile
xi2043 net8536 net8325 net8533 net8529 net8523 net8530 net8324 net8524 vdd vss unit_coupling_tile
xi2042 net8532 net8334 net8534 net8533 net8530 net8535 net8322 net8531 vdd vss unit_coupling_tile
xi2041 net8541 net8330 net8542 net8534 net8535 net8537 net8329 net8540 vdd vss unit_coupling_tile
xi2040 net8539 net8339 net8470 net8542 net8537 net8467 net8338 net8538 vdd vss unit_coupling_tile
xi2039 net8469 net8337 net8466 net8470 net8467 net8463 net8336 net8468 vdd vss unit_coupling_tile
xi2038 net8465 net8265 net8476 net8466 net8463 net8473 net8264 net8464 vdd vss unit_coupling_tile
xi2037 net8475 net8261 net8477 net8476 net8473 net8471 net8260 net8474 vdd vss unit_coupling_tile
xi2036 net8484 net8271 net8481 net8477 net8471 net8478 net8270 net8472 vdd vss unit_coupling_tile
xi2035 net8480 net8280 net8482 net8481 net8478 net8483 net8268 net8479 vdd vss unit_coupling_tile
xi2034 net8489 net8276 net8490 net8482 net8483 net8485 net8275 net8488 vdd vss unit_coupling_tile
xi2033 net8487 net8285 net8494 net8490 net8485 net8491 net8284 net8486 vdd vss unit_coupling_tile
xi2032 net8493 net8283 net8495 net8494 net8491 net8496 net8282 net8492 vdd vss unit_coupling_tile
xi2031 net8502 net8289 net8500 net8495 net8496 net8497 net8288 net8501 vdd vss unit_coupling_tile
xi2030 net8499 net8298 net8429 net8500 net8497 net8503 net8297 net8498 vdd vss unit_coupling_tile
xi2029 net8428 net8295 net8425 net8429 net8503 net8422 net8294 net8504 vdd vss unit_coupling_tile
xi2028 net8424 net8224 net8426 net8425 net8422 net8427 net8300 net8423 vdd vss unit_coupling_tile
xi2027 net8434 net8220 net8435 net8426 net8427 net8430 net8219 net8433 vdd vss unit_coupling_tile
xi2026 net8432 net8230 net8439 net8435 net8430 net8436 net8229 net8431 vdd vss unit_coupling_tile
xi2025 net8438 net8228 net8440 net8439 net8436 net8441 net8227 net8437 vdd vss unit_coupling_tile
xi2024 net8447 net8234 net8445 net8440 net8441 net8442 net8233 net8446 vdd vss unit_coupling_tile
xi2023 net8444 net8243 net8453 net8445 net8442 net8450 net8242 net8443 vdd vss unit_coupling_tile
xi2022 net8452 net8240 net8454 net8453 net8450 net8448 net8239 net8451 vdd vss unit_coupling_tile
xi2021 net8460 net8248 net8458 net8454 net8448 net8455 net8247 net8449 vdd vss unit_coupling_tile
xi2020 net8457 net8256 net8387 net8458 net8455 net8459 net8245 net8456 vdd vss unit_coupling_tile
xi2019 net8462 net8253 net8384 net8387 net8459 net8381 net8252 net8461 vdd vss unit_coupling_tile
xi2018 net8383 net8258 net8385 net8384 net8381 net8386 net8257 net8382 vdd vss unit_coupling_tile
xi2017 net8393 net8179 net8391 net8385 net8386 net8388 net8178 net8392 vdd vss unit_coupling_tile
xi2016 net8390 net8189 net8399 net8391 net8388 net8396 net8188 net8389 vdd vss unit_coupling_tile
xi2015 net8398 net8186 net8400 net8399 net8396 net8394 net8185 net8397 vdd vss unit_coupling_tile
xi2014 net8407 net8194 net8404 net8400 net8394 net8401 net8193 net8395 vdd vss unit_coupling_tile
xi2013 net8403 net8203 net8405 net8404 net8401 net8406 net8191 net8402 vdd vss unit_coupling_tile
xi2012 net8412 net8199 net8413 net8405 net8406 net8408 net8198 net8411 vdd vss unit_coupling_tile
xi2011 net8410 net8205 net8417 net8413 net8408 net8414 net8204 net8409 vdd vss unit_coupling_tile
xi2010 net8416 net8209 net8418 net8417 net8414 net8419 net8208 net8415 vdd vss unit_coupling_tile
xi2008 net8345 net8217 net8347 net8346 net8343 net8341 net8216 net8344 vdd vss unit_coupling_tile
xi2007 net8354 net8141 net8351 net8347 net8341 net8348 net8140 net8342 vdd vss unit_coupling_tile
xi2006 net8350 net8150 net8352 net8351 net8348 net8353 net8138 net8349 vdd vss unit_coupling_tile
xi2005 net8359 net8146 net8360 net8352 net8353 net8355 net8145 net8358 vdd vss unit_coupling_tile
xi2004 net8357 net8155 net8364 net8360 net8355 net8361 net8154 net8356 vdd vss unit_coupling_tile
xi2003 net8363 net8153 net8365 net8364 net8361 net8366 net8152 net8362 vdd vss unit_coupling_tile
xi2002 net8372 net8159 net8370 net8365 net8366 net8367 net8158 net8371 vdd vss unit_coupling_tile
xi2001 net8369 net8168 net8377 net8370 net8367 net8374 net8167 net8368 vdd vss unit_coupling_tile
xi2000 net8376 net8165 net8378 net8377 net8374 net8379 net8164 net8375 vdd vss unit_coupling_tile
xi1999 net8380 net8172 net8307 net63 net63 net8304 net8171 net8373 vdd vss unit_coupling_tile
xi1998 net8306 net8176 net8308 net8307 net8304 net8301 net8170 net8305 vdd vss unit_coupling_tile
xi1997 net8303 net8102 net8312 net8308 net8301 net8309 net8101 net8302 vdd vss unit_coupling_tile
xi1996 net8311 net8099 net8313 net8312 net8309 net8314 net8098 net8310 vdd vss unit_coupling_tile
xi1995 net8320 net8107 net8318 net8313 net8314 net8315 net8106 net8319 vdd vss unit_coupling_tile
xi1994 net8317 net8116 net8326 net8318 net8315 net8323 net8115 net8316 vdd vss unit_coupling_tile
xi1993 net8325 net8113 net8327 net8326 net8323 net8321 net8112 net8324 vdd vss unit_coupling_tile
xi1992 net8334 net8121 net8331 net8327 net8321 net8328 net8120 net8322 vdd vss unit_coupling_tile
xi1991 net8330 net8130 net8332 net8331 net8328 net8333 net8118 net8329 vdd vss unit_coupling_tile
xi1990 net8339 net8126 net8340 net8332 net8333 net8335 net8125 net8338 vdd vss unit_coupling_tile
xi1989 net8337 net8135 net8266 net8340 net8335 net8263 net8134 net8336 vdd vss unit_coupling_tile
xi1988 net8265 net8133 net8262 net8266 net8263 net8259 net8132 net8264 vdd vss unit_coupling_tile
xi1987 net8261 net8061 net8272 net8262 net8259 net8269 net8060 net8260 vdd vss unit_coupling_tile
xi1986 net8271 net8057 net8273 net8272 net8269 net8267 net8056 net8270 vdd vss unit_coupling_tile
xi1985 net8280 net8067 net8277 net8273 net8267 net8274 net8066 net8268 vdd vss unit_coupling_tile
xi1984 net8276 net8076 net8278 net8277 net8274 net8279 net8064 net8275 vdd vss unit_coupling_tile
xi1983 net8285 net8072 net8286 net8278 net8279 net8281 net8071 net8284 vdd vss unit_coupling_tile
xi1982 net8283 net8081 net8290 net8286 net8281 net8287 net8080 net8282 vdd vss unit_coupling_tile
xi1981 net8289 net8079 net8291 net8290 net8287 net8292 net8078 net8288 vdd vss unit_coupling_tile
xi1980 net8298 net8085 net8296 net8291 net8292 net8293 net8084 net8297 vdd vss unit_coupling_tile
xi1979 net8295 net8094 net8225 net8296 net8293 net8299 net8093 net8294 vdd vss unit_coupling_tile
xi1978 net8224 net8091 net8221 net8225 net8299 net8218 net8090 net8300 vdd vss unit_coupling_tile
xi1977 net8220 net8020 net8222 net8221 net8218 net8223 net8096 net8219 vdd vss unit_coupling_tile
xi1976 net8230 net8016 net8231 net8222 net8223 net8226 net8015 net8229 vdd vss unit_coupling_tile
xi1975 net8228 net8026 net8235 net8231 net8226 net8232 net8025 net8227 vdd vss unit_coupling_tile
xi1974 net8234 net8024 net8236 net8235 net8232 net8237 net8023 net8233 vdd vss unit_coupling_tile
xi1973 net8243 net8030 net8241 net8236 net8237 net8238 net8029 net8242 vdd vss unit_coupling_tile
xi1972 net8240 net8039 net8249 net8241 net8238 net8246 net8038 net8239 vdd vss unit_coupling_tile
xi1971 net8248 net8036 net8250 net8249 net8246 net8244 net8035 net8247 vdd vss unit_coupling_tile
xi1970 net8256 net8044 net8254 net8250 net8244 net8251 net8043 net8245 vdd vss unit_coupling_tile
xi1969 net8253 net8052 net8183 net8254 net8251 net8255 net8041 net8252 vdd vss unit_coupling_tile
xi1968 net8258 net8049 net8180 net8183 net8255 net8177 net8048 net8257 vdd vss unit_coupling_tile
xi1967 net8179 net8054 net8181 net8180 net8177 net8182 net8053 net8178 vdd vss unit_coupling_tile
xi1966 net8189 net7975 net8187 net8181 net8182 net8184 net7974 net8188 vdd vss unit_coupling_tile
xi1965 net8186 net7985 net8195 net8187 net8184 net8192 net7984 net8185 vdd vss unit_coupling_tile
xi1964 net8194 net7982 net8196 net8195 net8192 net8190 net7981 net8193 vdd vss unit_coupling_tile
xi1963 net8203 net7990 net8200 net8196 net8190 net8197 net7989 net8191 vdd vss unit_coupling_tile
xi1962 net8199 net7993 net8201 net8200 net8197 net8202 net7987 net8198 vdd vss unit_coupling_tile
xi1961 net8205 net7997 net8206 net8201 net8202 net8207 net7996 net8204 vdd vss unit_coupling_tile
xi1959 net8212 net8002 net8214 net8213 net8210 net8215 net8001 net8211 vdd vss unit_coupling_tile
xi1958 net8217 net8008 net8142 net8214 net8215 net8139 net8007 net8216 vdd vss unit_coupling_tile
xi1957 net8141 net8013 net8143 net8142 net8139 net8137 net8012 net8140 vdd vss unit_coupling_tile
xi1956 net8150 net7937 net8147 net8143 net8137 net8144 net7936 net8138 vdd vss unit_coupling_tile
xi1955 net8146 net7946 net8148 net8147 net8144 net8149 net7934 net8145 vdd vss unit_coupling_tile
xi1954 net8155 net7942 net8156 net8148 net8149 net8151 net7941 net8154 vdd vss unit_coupling_tile
xi1953 net8153 net7951 net8160 net8156 net8151 net8157 net7950 net8152 vdd vss unit_coupling_tile
xi1952 net8159 net7949 net8161 net8160 net8157 net8162 net7948 net8158 vdd vss unit_coupling_tile
xi1951 net8168 net7955 net8166 net8161 net8162 net8163 net7954 net8167 vdd vss unit_coupling_tile
xi1950 net8165 net7962 net8174 net8166 net8163 net8175 net7961 net8164 vdd vss unit_coupling_tile
xi1949 net8172 net7960 net8173 net64 net64 net8169 net7959 net8171 vdd vss unit_coupling_tile
xi1948 net8176 net7969 net8103 net8173 net8169 net8100 net7968 net8170 vdd vss unit_coupling_tile
xi1947 net8102 net7972 net8104 net8103 net8100 net8097 net7966 net8101 vdd vss unit_coupling_tile
xi1946 net8099 net7898 net8108 net8104 net8097 net8105 net7897 net8098 vdd vss unit_coupling_tile
xi1945 net8107 net7895 net8109 net8108 net8105 net8110 net7894 net8106 vdd vss unit_coupling_tile
xi1944 net8116 net7903 net8114 net8109 net8110 net8111 net7902 net8115 vdd vss unit_coupling_tile
xi1943 net8113 net7912 net8122 net8114 net8111 net8119 net7911 net8112 vdd vss unit_coupling_tile
xi1942 net8121 net7909 net8123 net8122 net8119 net8117 net7908 net8120 vdd vss unit_coupling_tile
xi1941 net8130 net7917 net8127 net8123 net8117 net8124 net7916 net8118 vdd vss unit_coupling_tile
xi1940 net8126 net7926 net8128 net8127 net8124 net8129 net7914 net8125 vdd vss unit_coupling_tile
xi1939 net8135 net7922 net8136 net8128 net8129 net8131 net7921 net8134 vdd vss unit_coupling_tile
xi1938 net8133 net7931 net8062 net8136 net8131 net8059 net7930 net8132 vdd vss unit_coupling_tile
xi1937 net8061 net7929 net8058 net8062 net8059 net8055 net7928 net8060 vdd vss unit_coupling_tile
xi1936 net8057 net7857 net8068 net8058 net8055 net8065 net7856 net8056 vdd vss unit_coupling_tile
xi1935 net8067 net7853 net8069 net8068 net8065 net8063 net7852 net8066 vdd vss unit_coupling_tile
xi1934 net8076 net7863 net8073 net8069 net8063 net8070 net7862 net8064 vdd vss unit_coupling_tile
xi1933 net8072 net7872 net8074 net8073 net8070 net8075 net7860 net8071 vdd vss unit_coupling_tile
xi1932 net8081 net7868 net8082 net8074 net8075 net8077 net7867 net8080 vdd vss unit_coupling_tile
xi1931 net8079 net7877 net8086 net8082 net8077 net8083 net7876 net8078 vdd vss unit_coupling_tile
xi1930 net8085 net7875 net8087 net8086 net8083 net8088 net7874 net8084 vdd vss unit_coupling_tile
xi1929 net8094 net7881 net8092 net8087 net8088 net8089 net7880 net8093 vdd vss unit_coupling_tile
xi1928 net8091 net7890 net8021 net8092 net8089 net8095 net7889 net8090 vdd vss unit_coupling_tile
xi1927 net8020 net7887 net8017 net8021 net8095 net8014 net7886 net8096 vdd vss unit_coupling_tile
xi1926 net8016 net7816 net8018 net8017 net8014 net8019 net7892 net8015 vdd vss unit_coupling_tile
xi1925 net8026 net7812 net8027 net8018 net8019 net8022 net7811 net8025 vdd vss unit_coupling_tile
xi1924 net8024 net7822 net8031 net8027 net8022 net8028 net7821 net8023 vdd vss unit_coupling_tile
xi1923 net8030 net7820 net8032 net8031 net8028 net8033 net7819 net8029 vdd vss unit_coupling_tile
xi1922 net8039 net7826 net8037 net8032 net8033 net8034 net7825 net8038 vdd vss unit_coupling_tile
xi1921 net8036 net7835 net8045 net8037 net8034 net8042 net7834 net8035 vdd vss unit_coupling_tile
xi1920 net8044 net7832 net8046 net8045 net8042 net8040 net7831 net8043 vdd vss unit_coupling_tile
xi1919 net8052 net7840 net8050 net8046 net8040 net8047 net7839 net8041 vdd vss unit_coupling_tile
xi1918 net8049 net7848 net7979 net8050 net8047 net8051 net7837 net8048 vdd vss unit_coupling_tile
xi1917 net8054 net7845 net7976 net7979 net8051 net7973 net7844 net8053 vdd vss unit_coupling_tile
xi1916 net7975 net7850 net7977 net7976 net7973 net7978 net7849 net7974 vdd vss unit_coupling_tile
xi1915 net7985 net7771 net7983 net7977 net7978 net7980 net7770 net7984 vdd vss unit_coupling_tile
xi1914 net7982 net7781 net7991 net7983 net7980 net7988 net7780 net7981 vdd vss unit_coupling_tile
xi1913 net7990 net7778 net7992 net7991 net7988 net7986 net7777 net7989 vdd vss unit_coupling_tile
xi1912 net7993 net7787 net7994 net7992 net7986 net7995 net7786 net7987 vdd vss unit_coupling_tile
xi1910 net8004 net7791 net8005 net7998 net7999 net8000 net7790 net8003 vdd vss unit_coupling_tile
xi1909 net8002 net7800 net8009 net8005 net8000 net8006 net7799 net8001 vdd vss unit_coupling_tile
xi1908 net8008 net7798 net8010 net8009 net8006 net8011 net7797 net8007 vdd vss unit_coupling_tile
xi1907 net8013 net7804 net7938 net8010 net8011 net7935 net7803 net8012 vdd vss unit_coupling_tile
xi1906 net7937 net7809 net7939 net7938 net7935 net7933 net7808 net7936 vdd vss unit_coupling_tile
xi1905 net7946 net7733 net7943 net7939 net7933 net7940 net7732 net7934 vdd vss unit_coupling_tile
xi1904 net7942 net7742 net7944 net7943 net7940 net7945 net7730 net7941 vdd vss unit_coupling_tile
xi1903 net7951 net7738 net7952 net7944 net7945 net7947 net7737 net7950 vdd vss unit_coupling_tile
xi1902 net7949 net7747 net7956 net7952 net7947 net7953 net7746 net7948 vdd vss unit_coupling_tile
xi1901 net7955 net7745 net7957 net7956 net7953 net7958 net7744 net7954 vdd vss unit_coupling_tile
xi1900 net7962 net7751 net7963 net7957 net7958 net7964 net7750 net7961 vdd vss unit_coupling_tile
xi1899 net7960 net7760 net7970 net65 net65 net7967 net7759 net7959 vdd vss unit_coupling_tile
xi1898 net7969 net7757 net7971 net7970 net7967 net7965 net7756 net7968 vdd vss unit_coupling_tile
xi1897 net7972 net7765 net7899 net7971 net7965 net7896 net7764 net7966 vdd vss unit_coupling_tile
xi1896 net7898 net7768 net7900 net7899 net7896 net7893 net7762 net7897 vdd vss unit_coupling_tile
xi1895 net7895 net7694 net7904 net7900 net7893 net7901 net7693 net7894 vdd vss unit_coupling_tile
xi1894 net7903 net7691 net7905 net7904 net7901 net7906 net7690 net7902 vdd vss unit_coupling_tile
xi1893 net7912 net7699 net7910 net7905 net7906 net7907 net7698 net7911 vdd vss unit_coupling_tile
xi1892 net7909 net7708 net7918 net7910 net7907 net7915 net7707 net7908 vdd vss unit_coupling_tile
xi1891 net7917 net7705 net7919 net7918 net7915 net7913 net7704 net7916 vdd vss unit_coupling_tile
xi1890 net7926 net7713 net7923 net7919 net7913 net7920 net7712 net7914 vdd vss unit_coupling_tile
xi1889 net7922 net7722 net7924 net7923 net7920 net7925 net7710 net7921 vdd vss unit_coupling_tile
xi1888 net7931 net7718 net7932 net7924 net7925 net7927 net7717 net7930 vdd vss unit_coupling_tile
xi1887 net7929 net7727 net7858 net7932 net7927 net7855 net7726 net7928 vdd vss unit_coupling_tile
xi1886 net7857 net7725 net7854 net7858 net7855 net7851 net7724 net7856 vdd vss unit_coupling_tile
xi1885 net7853 net7653 net7864 net7854 net7851 net7861 net7652 net7852 vdd vss unit_coupling_tile
xi1884 net7863 net7649 net7865 net7864 net7861 net7859 net7648 net7862 vdd vss unit_coupling_tile
xi1883 net7872 net7659 net7869 net7865 net7859 net7866 net7658 net7860 vdd vss unit_coupling_tile
xi1882 net7868 net7668 net7870 net7869 net7866 net7871 net7656 net7867 vdd vss unit_coupling_tile
xi1881 net7877 net7664 net7878 net7870 net7871 net7873 net7663 net7876 vdd vss unit_coupling_tile
xi1880 net7875 net7673 net7882 net7878 net7873 net7879 net7672 net7874 vdd vss unit_coupling_tile
xi1879 net7881 net7671 net7883 net7882 net7879 net7884 net7670 net7880 vdd vss unit_coupling_tile
xi1878 net7890 net7677 net7888 net7883 net7884 net7885 net7676 net7889 vdd vss unit_coupling_tile
xi1877 net7887 net7686 net7817 net7888 net7885 net7891 net7685 net7886 vdd vss unit_coupling_tile
xi1876 net7816 net7683 net7813 net7817 net7891 net7810 net7682 net7892 vdd vss unit_coupling_tile
xi1875 net7812 net7612 net7814 net7813 net7810 net7815 net7688 net7811 vdd vss unit_coupling_tile
xi1874 net7822 net7608 net7823 net7814 net7815 net7818 net7607 net7821 vdd vss unit_coupling_tile
xi1873 net7820 net7618 net7827 net7823 net7818 net7824 net7617 net7819 vdd vss unit_coupling_tile
xi1872 net7826 net7616 net7828 net7827 net7824 net7829 net7615 net7825 vdd vss unit_coupling_tile
xi1871 net7835 net7622 net7833 net7828 net7829 net7830 net7621 net7834 vdd vss unit_coupling_tile
xi1870 net7832 net7631 net7841 net7833 net7830 net7838 net7630 net7831 vdd vss unit_coupling_tile
xi1869 net7840 net7628 net7842 net7841 net7838 net7836 net7627 net7839 vdd vss unit_coupling_tile
xi1868 net7848 net7636 net7846 net7842 net7836 net7843 net7635 net7837 vdd vss unit_coupling_tile
xi1867 net7845 net7644 net7775 net7846 net7843 net7847 net7633 net7844 vdd vss unit_coupling_tile
xi1866 net7850 net7641 net7772 net7775 net7847 net7769 net7640 net7849 vdd vss unit_coupling_tile
xi1865 net7771 net7646 net7773 net7772 net7769 net7774 net7645 net7770 vdd vss unit_coupling_tile
xi1864 net7781 net7567 net7779 net7773 net7774 net7776 net7566 net7780 vdd vss unit_coupling_tile
xi1863 net7778 net7577 net7784 net7779 net7776 net7785 net7576 net7777 vdd vss unit_coupling_tile
xi1861 net7795 net7582 net7792 net7788 net7782 net7789 net7581 net7783 vdd vss unit_coupling_tile
xi1860 net7791 net7591 net7793 net7792 net7789 net7794 net7579 net7790 vdd vss unit_coupling_tile
xi1859 net7800 net7587 net7801 net7793 net7794 net7796 net7586 net7799 vdd vss unit_coupling_tile
xi1858 net7798 net7596 net7805 net7801 net7796 net7802 net7595 net7797 vdd vss unit_coupling_tile
xi1857 net7804 net7594 net7806 net7805 net7802 net7807 net7593 net7803 vdd vss unit_coupling_tile
xi1856 net7809 net7600 net7734 net7806 net7807 net7731 net7599 net7808 vdd vss unit_coupling_tile
xi1855 net7733 net7605 net7735 net7734 net7731 net7729 net7604 net7732 vdd vss unit_coupling_tile
xi1854 net7742 net7529 net7739 net7735 net7729 net7736 net7528 net7730 vdd vss unit_coupling_tile
xi1853 net7738 net7538 net7740 net7739 net7736 net7741 net7526 net7737 vdd vss unit_coupling_tile
xi1852 net7747 net7534 net7748 net7740 net7741 net7743 net7533 net7746 vdd vss unit_coupling_tile
xi1851 net7745 net7543 net7752 net7748 net7743 net7749 net7542 net7744 vdd vss unit_coupling_tile
xi1850 net7751 net7541 net7753 net7752 net7749 net7754 net7540 net7750 vdd vss unit_coupling_tile
xi1849 net7760 net7546 net7758 net66 net66 net7755 net7545 net7759 vdd vss unit_coupling_tile
xi1848 net7757 net7556 net7766 net7758 net7755 net7763 net7555 net7756 vdd vss unit_coupling_tile
xi1847 net7765 net7553 net7767 net7766 net7763 net7761 net7552 net7764 vdd vss unit_coupling_tile
xi1846 net7768 net7561 net7695 net7767 net7761 net7692 net7560 net7762 vdd vss unit_coupling_tile
xi1845 net7694 net7564 net7696 net7695 net7692 net7689 net7558 net7693 vdd vss unit_coupling_tile
xi1844 net7691 net7490 net7700 net7696 net7689 net7697 net7489 net7690 vdd vss unit_coupling_tile
xi1843 net7699 net7487 net7701 net7700 net7697 net7702 net7486 net7698 vdd vss unit_coupling_tile
xi1842 net7708 net7495 net7706 net7701 net7702 net7703 net7494 net7707 vdd vss unit_coupling_tile
xi1841 net7705 net7504 net7714 net7706 net7703 net7711 net7503 net7704 vdd vss unit_coupling_tile
xi1840 net7713 net7501 net7715 net7714 net7711 net7709 net7500 net7712 vdd vss unit_coupling_tile
xi1839 net7722 net7509 net7719 net7715 net7709 net7716 net7508 net7710 vdd vss unit_coupling_tile
xi1838 net7718 net7518 net7720 net7719 net7716 net7721 net7506 net7717 vdd vss unit_coupling_tile
xi1837 net7727 net7514 net7728 net7720 net7721 net7723 net7513 net7726 vdd vss unit_coupling_tile
xi1836 net7725 net7523 net7654 net7728 net7723 net7651 net7522 net7724 vdd vss unit_coupling_tile
xi1835 net7653 net7521 net7650 net7654 net7651 net7647 net7520 net7652 vdd vss unit_coupling_tile
xi1834 net7649 net7449 net7660 net7650 net7647 net7657 net7448 net7648 vdd vss unit_coupling_tile
xi1833 net7659 net7445 net7661 net7660 net7657 net7655 net7444 net7658 vdd vss unit_coupling_tile
xi1832 net7668 net7455 net7665 net7661 net7655 net7662 net7454 net7656 vdd vss unit_coupling_tile
xi1831 net7664 net7464 net7666 net7665 net7662 net7667 net7452 net7663 vdd vss unit_coupling_tile
xi1830 net7673 net7460 net7674 net7666 net7667 net7669 net7459 net7672 vdd vss unit_coupling_tile
xi1829 net7671 net7469 net7678 net7674 net7669 net7675 net7468 net7670 vdd vss unit_coupling_tile
xi1828 net7677 net7467 net7679 net7678 net7675 net7680 net7466 net7676 vdd vss unit_coupling_tile
xi1827 net7686 net7473 net7684 net7679 net7680 net7681 net7472 net7685 vdd vss unit_coupling_tile
xi1826 net7683 net7482 net7613 net7684 net7681 net7687 net7481 net7682 vdd vss unit_coupling_tile
xi1825 net7612 net7479 net7609 net7613 net7687 net7606 net7478 net7688 vdd vss unit_coupling_tile
xi1824 net7608 net7408 net7610 net7609 net7606 net7611 net7484 net7607 vdd vss unit_coupling_tile
xi1823 net7618 net7404 net7619 net7610 net7611 net7614 net7403 net7617 vdd vss unit_coupling_tile
xi1822 net7616 net7414 net7623 net7619 net7614 net7620 net7413 net7615 vdd vss unit_coupling_tile
xi1821 net7622 net7412 net7624 net7623 net7620 net7625 net7411 net7621 vdd vss unit_coupling_tile
xi1820 net7631 net7418 net7629 net7624 net7625 net7626 net7417 net7630 vdd vss unit_coupling_tile
xi1819 net7628 net7427 net7637 net7629 net7626 net7634 net7426 net7627 vdd vss unit_coupling_tile
xi1818 net7636 net7424 net7638 net7637 net7634 net7632 net7423 net7635 vdd vss unit_coupling_tile
xi1817 net7644 net7432 net7642 net7638 net7632 net7639 net7431 net7633 vdd vss unit_coupling_tile
xi1816 net7641 net7440 net7571 net7642 net7639 net7643 net7429 net7640 vdd vss unit_coupling_tile
xi1815 net7646 net7437 net7568 net7571 net7643 net7565 net7436 net7645 vdd vss unit_coupling_tile
xi1814 net7567 net7442 net7569 net7568 net7565 net7570 net7441 net7566 vdd vss unit_coupling_tile
xi1812 net7574 net7373 net7583 net7575 net7572 net7580 net7372 net7573 vdd vss unit_coupling_tile
xi1811 net7582 net7370 net7584 net7583 net7580 net7578 net7369 net7581 vdd vss unit_coupling_tile
xi1810 net7591 net7378 net7588 net7584 net7578 net7585 net7377 net7579 vdd vss unit_coupling_tile
xi1809 net7587 net7387 net7589 net7588 net7585 net7590 net7375 net7586 vdd vss unit_coupling_tile
xi1808 net7596 net7383 net7597 net7589 net7590 net7592 net7382 net7595 vdd vss unit_coupling_tile
xi1807 net7594 net7392 net7601 net7597 net7592 net7598 net7391 net7593 vdd vss unit_coupling_tile
xi1806 net7600 net7390 net7602 net7601 net7598 net7603 net7389 net7599 vdd vss unit_coupling_tile
xi1805 net7605 net7396 net7530 net7602 net7603 net7527 net7395 net7604 vdd vss unit_coupling_tile
xi1804 net7529 net7401 net7531 net7530 net7527 net7525 net7400 net7528 vdd vss unit_coupling_tile
xi1803 net7538 net7325 net7535 net7531 net7525 net7532 net7324 net7526 vdd vss unit_coupling_tile
xi1802 net7534 net7334 net7536 net7535 net7532 net7537 net7322 net7533 vdd vss unit_coupling_tile
xi1801 net7543 net7330 net7544 net7536 net7537 net7539 net7329 net7542 vdd vss unit_coupling_tile
xi1800 net7541 net7338 net7549 net7544 net7539 net7550 net7337 net7540 vdd vss unit_coupling_tile
xi1799 net7546 net7336 net7547 net67 net67 net7548 net7335 net7545 vdd vss unit_coupling_tile
xi1798 net7556 net7343 net7554 net7547 net7548 net7551 net7342 net7555 vdd vss unit_coupling_tile
xi1797 net7553 net7352 net7562 net7554 net7551 net7559 net7351 net7552 vdd vss unit_coupling_tile
xi1796 net7561 net7349 net7563 net7562 net7559 net7557 net7348 net7560 vdd vss unit_coupling_tile
xi1795 net7564 net7357 net7491 net7563 net7557 net7488 net7356 net7558 vdd vss unit_coupling_tile
xi1794 net7490 net7360 net7492 net7491 net7488 net7485 net7354 net7489 vdd vss unit_coupling_tile
xi1793 net7487 net7286 net7496 net7492 net7485 net7493 net7285 net7486 vdd vss unit_coupling_tile
xi1792 net7495 net7283 net7497 net7496 net7493 net7498 net7282 net7494 vdd vss unit_coupling_tile
xi1791 net7504 net7291 net7502 net7497 net7498 net7499 net7290 net7503 vdd vss unit_coupling_tile
xi1790 net7501 net7300 net7510 net7502 net7499 net7507 net7299 net7500 vdd vss unit_coupling_tile
xi1789 net7509 net7297 net7511 net7510 net7507 net7505 net7296 net7508 vdd vss unit_coupling_tile
xi1788 net7518 net7305 net7515 net7511 net7505 net7512 net7304 net7506 vdd vss unit_coupling_tile
xi1787 net7514 net7314 net7516 net7515 net7512 net7517 net7302 net7513 vdd vss unit_coupling_tile
xi1786 net7523 net7310 net7524 net7516 net7517 net7519 net7309 net7522 vdd vss unit_coupling_tile
xi1785 net7521 net7319 net7450 net7524 net7519 net7447 net7318 net7520 vdd vss unit_coupling_tile
xi1784 net7449 net7317 net7446 net7450 net7447 net7443 net7316 net7448 vdd vss unit_coupling_tile
xi1783 net7445 net7245 net7456 net7446 net7443 net7453 net7244 net7444 vdd vss unit_coupling_tile
xi1782 net7455 net7241 net7457 net7456 net7453 net7451 net7240 net7454 vdd vss unit_coupling_tile
xi1781 net7464 net7251 net7461 net7457 net7451 net7458 net7250 net7452 vdd vss unit_coupling_tile
xi1780 net7460 net7260 net7462 net7461 net7458 net7463 net7248 net7459 vdd vss unit_coupling_tile
xi1779 net7469 net7256 net7470 net7462 net7463 net7465 net7255 net7468 vdd vss unit_coupling_tile
xi1778 net7467 net7265 net7474 net7470 net7465 net7471 net7264 net7466 vdd vss unit_coupling_tile
xi1777 net7473 net7263 net7475 net7474 net7471 net7476 net7262 net7472 vdd vss unit_coupling_tile
xi1776 net7482 net7269 net7480 net7475 net7476 net7477 net7268 net7481 vdd vss unit_coupling_tile
xi1775 net7479 net7278 net7409 net7480 net7477 net7483 net7277 net7478 vdd vss unit_coupling_tile
xi1774 net7408 net7275 net7405 net7409 net7483 net7402 net7274 net7484 vdd vss unit_coupling_tile
xi1773 net7404 net7204 net7406 net7405 net7402 net7407 net7280 net7403 vdd vss unit_coupling_tile
xi1772 net7414 net7200 net7415 net7406 net7407 net7410 net7199 net7413 vdd vss unit_coupling_tile
xi1771 net7412 net7210 net7419 net7415 net7410 net7416 net7209 net7411 vdd vss unit_coupling_tile
xi1770 net7418 net7208 net7420 net7419 net7416 net7421 net7207 net7417 vdd vss unit_coupling_tile
xi1769 net7427 net7214 net7425 net7420 net7421 net7422 net7213 net7426 vdd vss unit_coupling_tile
xi1768 net7424 net7223 net7433 net7425 net7422 net7430 net7222 net7423 vdd vss unit_coupling_tile
xi1767 net7432 net7220 net7434 net7433 net7430 net7428 net7219 net7431 vdd vss unit_coupling_tile
xi1766 net7440 net7226 net7438 net7434 net7428 net7435 net7225 net7429 vdd vss unit_coupling_tile
xi1765 net7437 net7236 net7367 net7438 net7435 net7439 net7230 net7436 vdd vss unit_coupling_tile
xi1763 net7363 net7238 net7365 net7364 net7361 net7366 net7237 net7362 vdd vss unit_coupling_tile
xi1762 net7373 net7159 net7371 net7365 net7366 net7368 net7158 net7372 vdd vss unit_coupling_tile
xi1761 net7370 net7169 net7379 net7371 net7368 net7376 net7168 net7369 vdd vss unit_coupling_tile
xi1760 net7378 net7166 net7380 net7379 net7376 net7374 net7165 net7377 vdd vss unit_coupling_tile
xi1759 net7387 net7174 net7384 net7380 net7374 net7381 net7173 net7375 vdd vss unit_coupling_tile
xi1758 net7383 net7183 net7385 net7384 net7381 net7386 net7171 net7382 vdd vss unit_coupling_tile
xi1757 net7392 net7179 net7393 net7385 net7386 net7388 net7178 net7391 vdd vss unit_coupling_tile
xi1756 net7390 net7188 net7397 net7393 net7388 net7394 net7187 net7389 vdd vss unit_coupling_tile
xi1755 net7396 net7186 net7398 net7397 net7394 net7399 net7185 net7395 vdd vss unit_coupling_tile
xi1754 net7401 net7192 net7326 net7398 net7399 net7323 net7191 net7400 vdd vss unit_coupling_tile
xi1753 net7325 net7197 net7327 net7326 net7323 net7321 net7196 net7324 vdd vss unit_coupling_tile
xi1752 net7334 net7121 net7331 net7327 net7321 net7328 net7120 net7322 vdd vss unit_coupling_tile
xi1751 net7330 net7130 net7332 net7331 net7328 net7333 net7118 net7329 vdd vss unit_coupling_tile
xi1750 net7338 net7126 net7339 net7332 net7333 net7340 net7125 net7337 vdd vss unit_coupling_tile
xi1749 net7336 net7135 net7344 net68 net68 net7341 net7134 net7335 vdd vss unit_coupling_tile
xi1748 net7343 net7133 net7345 net7344 net7341 net7346 net7132 net7342 vdd vss unit_coupling_tile
xi1747 net7352 net7139 net7350 net7345 net7346 net7347 net7138 net7351 vdd vss unit_coupling_tile
xi1746 net7349 net7148 net7358 net7350 net7347 net7355 net7147 net7348 vdd vss unit_coupling_tile
xi1745 net7357 net7145 net7359 net7358 net7355 net7353 net7144 net7356 vdd vss unit_coupling_tile
xi1744 net7360 net7153 net7287 net7359 net7353 net7284 net7152 net7354 vdd vss unit_coupling_tile
xi1743 net7286 net7156 net7288 net7287 net7284 net7281 net7150 net7285 vdd vss unit_coupling_tile
xi1742 net7283 net7082 net7292 net7288 net7281 net7289 net7081 net7282 vdd vss unit_coupling_tile
xi1741 net7291 net7079 net7293 net7292 net7289 net7294 net7078 net7290 vdd vss unit_coupling_tile
xi1740 net7300 net7087 net7298 net7293 net7294 net7295 net7086 net7299 vdd vss unit_coupling_tile
xi1739 net7297 net7096 net7306 net7298 net7295 net7303 net7095 net7296 vdd vss unit_coupling_tile
xi1738 net7305 net7093 net7307 net7306 net7303 net7301 net7092 net7304 vdd vss unit_coupling_tile
xi1737 net7314 net7101 net7311 net7307 net7301 net7308 net7100 net7302 vdd vss unit_coupling_tile
xi1736 net7310 net7110 net7312 net7311 net7308 net7313 net7098 net7309 vdd vss unit_coupling_tile
xi1735 net7319 net7106 net7320 net7312 net7313 net7315 net7105 net7318 vdd vss unit_coupling_tile
xi1734 net7317 net7115 net7246 net7320 net7315 net7243 net7114 net7316 vdd vss unit_coupling_tile
xi1733 net7245 net7113 net7242 net7246 net7243 net7239 net7112 net7244 vdd vss unit_coupling_tile
xi1732 net7241 net7041 net7252 net7242 net7239 net7249 net7040 net7240 vdd vss unit_coupling_tile
xi1731 net7251 net7037 net7253 net7252 net7249 net7247 net7036 net7250 vdd vss unit_coupling_tile
xi1730 net7260 net7047 net7257 net7253 net7247 net7254 net7046 net7248 vdd vss unit_coupling_tile
xi1729 net7256 net7056 net7258 net7257 net7254 net7259 net7044 net7255 vdd vss unit_coupling_tile
xi1728 net7265 net7052 net7266 net7258 net7259 net7261 net7051 net7264 vdd vss unit_coupling_tile
xi1727 net7263 net7061 net7270 net7266 net7261 net7267 net7060 net7262 vdd vss unit_coupling_tile
xi1726 net7269 net7059 net7271 net7270 net7267 net7272 net7058 net7268 vdd vss unit_coupling_tile
xi1725 net7278 net7065 net7276 net7271 net7272 net7273 net7064 net7277 vdd vss unit_coupling_tile
xi1724 net7275 net7074 net7205 net7276 net7273 net7279 net7073 net7274 vdd vss unit_coupling_tile
xi1723 net7204 net7071 net7201 net7205 net7279 net7198 net7070 net7280 vdd vss unit_coupling_tile
xi1722 net7200 net7000 net7202 net7201 net7198 net7203 net7076 net7199 vdd vss unit_coupling_tile
xi1721 net7210 net6996 net7211 net7202 net7203 net7206 net6995 net7209 vdd vss unit_coupling_tile
xi1720 net7208 net7006 net7215 net7211 net7206 net7212 net7005 net7207 vdd vss unit_coupling_tile
xi1719 net7214 net7004 net7216 net7215 net7212 net7217 net7003 net7213 vdd vss unit_coupling_tile
xi1718 net7223 net7010 net7221 net7216 net7217 net7218 net7009 net7222 vdd vss unit_coupling_tile
xi1717 net7220 net7015 net7227 net7221 net7218 net7224 net7014 net7219 vdd vss unit_coupling_tile
xi1716 net7226 net7019 net7228 net7227 net7224 net7229 net7018 net7225 vdd vss unit_coupling_tile
xi1714 net7233 net7032 net7163 net7234 net7231 net7235 net7021 net7232 vdd vss unit_coupling_tile
xi1713 net7238 net7029 net7160 net7163 net7235 net7157 net7028 net7237 vdd vss unit_coupling_tile
xi1712 net7159 net7034 net7161 net7160 net7157 net7162 net7033 net7158 vdd vss unit_coupling_tile
xi1711 net7169 net6955 net7167 net7161 net7162 net7164 net6954 net7168 vdd vss unit_coupling_tile
xi1710 net7166 net6965 net7175 net7167 net7164 net7172 net6964 net7165 vdd vss unit_coupling_tile
xi1709 net7174 net6962 net7176 net7175 net7172 net7170 net6961 net7173 vdd vss unit_coupling_tile
xi1708 net7183 net6970 net7180 net7176 net7170 net7177 net6969 net7171 vdd vss unit_coupling_tile
xi1707 net7179 net6979 net7181 net7180 net7177 net7182 net6967 net7178 vdd vss unit_coupling_tile
xi1706 net7188 net6975 net7189 net7181 net7182 net7184 net6974 net7187 vdd vss unit_coupling_tile
xi1705 net7186 net6984 net7193 net7189 net7184 net7190 net6983 net7185 vdd vss unit_coupling_tile
xi1704 net7192 net6982 net7194 net7193 net7190 net7195 net6981 net7191 vdd vss unit_coupling_tile
xi1703 net7197 net6988 net7122 net7194 net7195 net7119 net6987 net7196 vdd vss unit_coupling_tile
xi1702 net7121 net6993 net7123 net7122 net7119 net7117 net6992 net7120 vdd vss unit_coupling_tile
xi1701 net7130 net6917 net7127 net7123 net7117 net7124 net6916 net7118 vdd vss unit_coupling_tile
xi1700 net7126 net6924 net7128 net7127 net7124 net7129 net6914 net7125 vdd vss unit_coupling_tile
xi1699 net7135 net6921 net7136 net69 net69 net7131 net6920 net7134 vdd vss unit_coupling_tile
xi1698 net7133 net6931 net7140 net7136 net7131 net7137 net6930 net7132 vdd vss unit_coupling_tile
xi1697 net7139 net6929 net7141 net7140 net7137 net7142 net6928 net7138 vdd vss unit_coupling_tile
xi1696 net7148 net6935 net7146 net7141 net7142 net7143 net6934 net7147 vdd vss unit_coupling_tile
xi1695 net7145 net6944 net7154 net7146 net7143 net7151 net6943 net7144 vdd vss unit_coupling_tile
xi1694 net7153 net6941 net7155 net7154 net7151 net7149 net6940 net7152 vdd vss unit_coupling_tile
xi1693 net7156 net6949 net7083 net7155 net7149 net7080 net6948 net7150 vdd vss unit_coupling_tile
xi1692 net7082 net6952 net7084 net7083 net7080 net7077 net6946 net7081 vdd vss unit_coupling_tile
xi1691 net7079 net6878 net7088 net7084 net7077 net7085 net6877 net7078 vdd vss unit_coupling_tile
xi1690 net7087 net6875 net7089 net7088 net7085 net7090 net6874 net7086 vdd vss unit_coupling_tile
xi1689 net7096 net6883 net7094 net7089 net7090 net7091 net6882 net7095 vdd vss unit_coupling_tile
xi1688 net7093 net6892 net7102 net7094 net7091 net7099 net6891 net7092 vdd vss unit_coupling_tile
xi1687 net7101 net6889 net7103 net7102 net7099 net7097 net6888 net7100 vdd vss unit_coupling_tile
xi1686 net7110 net6897 net7107 net7103 net7097 net7104 net6896 net7098 vdd vss unit_coupling_tile
xi1685 net7106 net6906 net7108 net7107 net7104 net7109 net6894 net7105 vdd vss unit_coupling_tile
xi1684 net7115 net6902 net7116 net7108 net7109 net7111 net6901 net7114 vdd vss unit_coupling_tile
xi1683 net7113 net6911 net7042 net7116 net7111 net7039 net6910 net7112 vdd vss unit_coupling_tile
xi1682 net7041 net6909 net7038 net7042 net7039 net7035 net6908 net7040 vdd vss unit_coupling_tile
xi1681 net7037 net6837 net7048 net7038 net7035 net7045 net6836 net7036 vdd vss unit_coupling_tile
xi1680 net7047 net6833 net7049 net7048 net7045 net7043 net6832 net7046 vdd vss unit_coupling_tile
xi1679 net7056 net6843 net7053 net7049 net7043 net7050 net6842 net7044 vdd vss unit_coupling_tile
xi1678 net7052 net6852 net7054 net7053 net7050 net7055 net6840 net7051 vdd vss unit_coupling_tile
xi1677 net7061 net6848 net7062 net7054 net7055 net7057 net6847 net7060 vdd vss unit_coupling_tile
xi1676 net7059 net6857 net7066 net7062 net7057 net7063 net6856 net7058 vdd vss unit_coupling_tile
xi1675 net7065 net6855 net7067 net7066 net7063 net7068 net6854 net7064 vdd vss unit_coupling_tile
xi1674 net7074 net6861 net7072 net7067 net7068 net7069 net6860 net7073 vdd vss unit_coupling_tile
xi1673 net7071 net6870 net7001 net7072 net7069 net7075 net6869 net7070 vdd vss unit_coupling_tile
xi1672 net7000 net6867 net6997 net7001 net7075 net6994 net6866 net7076 vdd vss unit_coupling_tile
xi1671 net6996 net6796 net6998 net6997 net6994 net6999 net6872 net6995 vdd vss unit_coupling_tile
xi1670 net7006 net6792 net7007 net6998 net6999 net7002 net6791 net7005 vdd vss unit_coupling_tile
xi1669 net7004 net6802 net7011 net7007 net7002 net7008 net6801 net7003 vdd vss unit_coupling_tile
xi1668 net7010 net6800 net7012 net7011 net7008 net7013 net6799 net7009 vdd vss unit_coupling_tile
xi1667 net7015 net6807 net7016 net7012 net7013 net7017 net6806 net7014 vdd vss unit_coupling_tile
xi1665 net7024 net6812 net7026 net7025 net7022 net7020 net6811 net7023 vdd vss unit_coupling_tile
xi1664 net7032 net6820 net7030 net7026 net7020 net7027 net6819 net7021 vdd vss unit_coupling_tile
xi1663 net7029 net6828 net6959 net7030 net7027 net7031 net6817 net7028 vdd vss unit_coupling_tile
xi1662 net7034 net6825 net6956 net6959 net7031 net6953 net6824 net7033 vdd vss unit_coupling_tile
xi1661 net6955 net6830 net6957 net6956 net6953 net6958 net6829 net6954 vdd vss unit_coupling_tile
xi1660 net6965 net6751 net6963 net6957 net6958 net6960 net6750 net6964 vdd vss unit_coupling_tile
xi1659 net6962 net6761 net6971 net6963 net6960 net6968 net6760 net6961 vdd vss unit_coupling_tile
xi1658 net6970 net6758 net6972 net6971 net6968 net6966 net6757 net6969 vdd vss unit_coupling_tile
xi1657 net6979 net6766 net6976 net6972 net6966 net6973 net6765 net6967 vdd vss unit_coupling_tile
xi1656 net6975 net6775 net6977 net6976 net6973 net6978 net6763 net6974 vdd vss unit_coupling_tile
xi1655 net6984 net6771 net6985 net6977 net6978 net6980 net6770 net6983 vdd vss unit_coupling_tile
xi1654 net6982 net6780 net6989 net6985 net6980 net6986 net6779 net6981 vdd vss unit_coupling_tile
xi1653 net6988 net6778 net6990 net6989 net6986 net6991 net6777 net6987 vdd vss unit_coupling_tile
xi1652 net6993 net6784 net6918 net6990 net6991 net6915 net6783 net6992 vdd vss unit_coupling_tile
xi1651 net6917 net6789 net6919 net6918 net6915 net6913 net6788 net6916 vdd vss unit_coupling_tile
xi1650 net6924 net6712 net6925 net6919 net6913 net6926 net6711 net6914 vdd vss unit_coupling_tile
xi1649 net6921 net6722 net6922 net70 net70 net6923 net6709 net6920 vdd vss unit_coupling_tile
xi1648 net6931 net6718 net6932 net6922 net6923 net6927 net6717 net6930 vdd vss unit_coupling_tile
xi1647 net6929 net6727 net6936 net6932 net6927 net6933 net6726 net6928 vdd vss unit_coupling_tile
xi1646 net6935 net6725 net6937 net6936 net6933 net6938 net6724 net6934 vdd vss unit_coupling_tile
xi1645 net6944 net6731 net6942 net6937 net6938 net6939 net6730 net6943 vdd vss unit_coupling_tile
xi1644 net6941 net6740 net6950 net6942 net6939 net6947 net6739 net6940 vdd vss unit_coupling_tile
xi1643 net6949 net6737 net6951 net6950 net6947 net6945 net6736 net6948 vdd vss unit_coupling_tile
xi1642 net6952 net6745 net6879 net6951 net6945 net6876 net6744 net6946 vdd vss unit_coupling_tile
xi1641 net6878 net6748 net6880 net6879 net6876 net6873 net6742 net6877 vdd vss unit_coupling_tile
xi1640 net6875 net6674 net6884 net6880 net6873 net6881 net6673 net6874 vdd vss unit_coupling_tile
xi1639 net6883 net6671 net6885 net6884 net6881 net6886 net6670 net6882 vdd vss unit_coupling_tile
xi1638 net6892 net6679 net6890 net6885 net6886 net6887 net6678 net6891 vdd vss unit_coupling_tile
xi1637 net6889 net6688 net6898 net6890 net6887 net6895 net6687 net6888 vdd vss unit_coupling_tile
xi1636 net6897 net6685 net6899 net6898 net6895 net6893 net6684 net6896 vdd vss unit_coupling_tile
xi1635 net6906 net6693 net6903 net6899 net6893 net6900 net6692 net6894 vdd vss unit_coupling_tile
xi1634 net6902 net6702 net6904 net6903 net6900 net6905 net6690 net6901 vdd vss unit_coupling_tile
xi1633 net6911 net6698 net6912 net6904 net6905 net6907 net6697 net6910 vdd vss unit_coupling_tile
xi1632 net6909 net6707 net6838 net6912 net6907 net6835 net6706 net6908 vdd vss unit_coupling_tile
xi1631 net6837 net6705 net6834 net6838 net6835 net6831 net6704 net6836 vdd vss unit_coupling_tile
xi1630 net6833 net6633 net6844 net6834 net6831 net6841 net6632 net6832 vdd vss unit_coupling_tile
xi1629 net6843 net6629 net6845 net6844 net6841 net6839 net6628 net6842 vdd vss unit_coupling_tile
xi1628 net6852 net6639 net6849 net6845 net6839 net6846 net6638 net6840 vdd vss unit_coupling_tile
xi1627 net6848 net6648 net6850 net6849 net6846 net6851 net6636 net6847 vdd vss unit_coupling_tile
xi1626 net6857 net6644 net6858 net6850 net6851 net6853 net6643 net6856 vdd vss unit_coupling_tile
xi1625 net6855 net6653 net6862 net6858 net6853 net6859 net6652 net6854 vdd vss unit_coupling_tile
xi1624 net6861 net6651 net6863 net6862 net6859 net6864 net6650 net6860 vdd vss unit_coupling_tile
xi1623 net6870 net6657 net6868 net6863 net6864 net6865 net6656 net6869 vdd vss unit_coupling_tile
xi1622 net6867 net6666 net6797 net6868 net6865 net6871 net6665 net6866 vdd vss unit_coupling_tile
xi1621 net6796 net6663 net6793 net6797 net6871 net6790 net6662 net6872 vdd vss unit_coupling_tile
xi1620 net6792 net6592 net6794 net6793 net6790 net6795 net6668 net6791 vdd vss unit_coupling_tile
xi1619 net6802 net6588 net6803 net6794 net6795 net6798 net6587 net6801 vdd vss unit_coupling_tile
xi1618 net6800 net6598 net6804 net6803 net6798 net6805 net6597 net6799 vdd vss unit_coupling_tile
xi1616 net6815 net6602 net6813 net6808 net6809 net6810 net6601 net6814 vdd vss unit_coupling_tile
xi1615 net6812 net6611 net6821 net6813 net6810 net6818 net6610 net6811 vdd vss unit_coupling_tile
xi1614 net6820 net6608 net6822 net6821 net6818 net6816 net6607 net6819 vdd vss unit_coupling_tile
xi1613 net6828 net6616 net6826 net6822 net6816 net6823 net6615 net6817 vdd vss unit_coupling_tile
xi1612 net6825 net6624 net6755 net6826 net6823 net6827 net6613 net6824 vdd vss unit_coupling_tile
xi1611 net6830 net6621 net6752 net6755 net6827 net6749 net6620 net6829 vdd vss unit_coupling_tile
xi1610 net6751 net6626 net6753 net6752 net6749 net6754 net6625 net6750 vdd vss unit_coupling_tile
xi1609 net6761 net6547 net6759 net6753 net6754 net6756 net6546 net6760 vdd vss unit_coupling_tile
xi1608 net6758 net6557 net6767 net6759 net6756 net6764 net6556 net6757 vdd vss unit_coupling_tile
xi1607 net6766 net6554 net6768 net6767 net6764 net6762 net6553 net6765 vdd vss unit_coupling_tile
xi1606 net6775 net6562 net6772 net6768 net6762 net6769 net6561 net6763 vdd vss unit_coupling_tile
xi1605 net6771 net6571 net6773 net6772 net6769 net6774 net6559 net6770 vdd vss unit_coupling_tile
xi1604 net6780 net6567 net6781 net6773 net6774 net6776 net6566 net6779 vdd vss unit_coupling_tile
xi1603 net6778 net6576 net6785 net6781 net6776 net6782 net6575 net6777 vdd vss unit_coupling_tile
xi1602 net6784 net6574 net6786 net6785 net6782 net6787 net6573 net6783 vdd vss unit_coupling_tile
xi1601 net6789 net6580 net6713 net6786 net6787 net6710 net6579 net6788 vdd vss unit_coupling_tile
xi1600 net6712 net6585 net6714 net6713 net6710 net6715 net6584 net6711 vdd vss unit_coupling_tile
xi1599 net6722 net6508 net6719 net71 net71 net6716 net6507 net6709 vdd vss unit_coupling_tile
xi1598 net6718 net6518 net6720 net6719 net6716 net6721 net6506 net6717 vdd vss unit_coupling_tile
xi1597 net6727 net6514 net6728 net6720 net6721 net6723 net6513 net6726 vdd vss unit_coupling_tile
xi1596 net6725 net6523 net6732 net6728 net6723 net6729 net6522 net6724 vdd vss unit_coupling_tile
xi1595 net6731 net6521 net6733 net6732 net6729 net6734 net6520 net6730 vdd vss unit_coupling_tile
xi1594 net6740 net6527 net6738 net6733 net6734 net6735 net6526 net6739 vdd vss unit_coupling_tile
xi1593 net6737 net6536 net6746 net6738 net6735 net6743 net6535 net6736 vdd vss unit_coupling_tile
xi1592 net6745 net6533 net6747 net6746 net6743 net6741 net6532 net6744 vdd vss unit_coupling_tile
xi1591 net6748 net6541 net6675 net6747 net6741 net6672 net6540 net6742 vdd vss unit_coupling_tile
xi1590 net6674 net6544 net6676 net6675 net6672 net6669 net6538 net6673 vdd vss unit_coupling_tile
xi1589 net6671 net6470 net6680 net6676 net6669 net6677 net6469 net6670 vdd vss unit_coupling_tile
xi1588 net6679 net6467 net6681 net6680 net6677 net6682 net6466 net6678 vdd vss unit_coupling_tile
xi1587 net6688 net6475 net6686 net6681 net6682 net6683 net6474 net6687 vdd vss unit_coupling_tile
xi1586 net6685 net6484 net6694 net6686 net6683 net6691 net6483 net6684 vdd vss unit_coupling_tile
xi1585 net6693 net6481 net6695 net6694 net6691 net6689 net6480 net6692 vdd vss unit_coupling_tile
xi1584 net6702 net6489 net6699 net6695 net6689 net6696 net6488 net6690 vdd vss unit_coupling_tile
xi1583 net6698 net6498 net6700 net6699 net6696 net6701 net6486 net6697 vdd vss unit_coupling_tile
xi1582 net6707 net6494 net6708 net6700 net6701 net6703 net6493 net6706 vdd vss unit_coupling_tile
xi1581 net6705 net6503 net6634 net6708 net6703 net6631 net6502 net6704 vdd vss unit_coupling_tile
xi1580 net6633 net6501 net6630 net6634 net6631 net6627 net6500 net6632 vdd vss unit_coupling_tile
xi1579 net6629 net6429 net6640 net6630 net6627 net6637 net6428 net6628 vdd vss unit_coupling_tile
xi1578 net6639 net6425 net6641 net6640 net6637 net6635 net6424 net6638 vdd vss unit_coupling_tile
xi1577 net6648 net6435 net6645 net6641 net6635 net6642 net6434 net6636 vdd vss unit_coupling_tile
xi1576 net6644 net6444 net6646 net6645 net6642 net6647 net6432 net6643 vdd vss unit_coupling_tile
xi1575 net6653 net6440 net6654 net6646 net6647 net6649 net6439 net6652 vdd vss unit_coupling_tile
xi1574 net6651 net6449 net6658 net6654 net6649 net6655 net6448 net6650 vdd vss unit_coupling_tile
xi1573 net6657 net6447 net6659 net6658 net6655 net6660 net6446 net6656 vdd vss unit_coupling_tile
xi1572 net6666 net6453 net6664 net6659 net6660 net6661 net6452 net6665 vdd vss unit_coupling_tile
xi1571 net6663 net6462 net6593 net6664 net6661 net6667 net6461 net6662 vdd vss unit_coupling_tile
xi1570 net6592 net6459 net6589 net6593 net6667 net6586 net6458 net6668 vdd vss unit_coupling_tile
xi1569 net6588 net6388 net6590 net6589 net6586 net6591 net6464 net6587 vdd vss unit_coupling_tile
xi1567 net6596 net6394 net6603 net6599 net6594 net6600 net6393 net6595 vdd vss unit_coupling_tile
xi1566 net6602 net6392 net6604 net6603 net6600 net6605 net6391 net6601 vdd vss unit_coupling_tile
xi1565 net6611 net6398 net6609 net6604 net6605 net6606 net6397 net6610 vdd vss unit_coupling_tile
xi1564 net6608 net6407 net6617 net6609 net6606 net6614 net6406 net6607 vdd vss unit_coupling_tile
xi1563 net6616 net6404 net6618 net6617 net6614 net6612 net6403 net6615 vdd vss unit_coupling_tile
xi1562 net6624 net6412 net6622 net6618 net6612 net6619 net6411 net6613 vdd vss unit_coupling_tile
xi1561 net6621 net6420 net6551 net6622 net6619 net6623 net6409 net6620 vdd vss unit_coupling_tile
xi1560 net6626 net6417 net6548 net6551 net6623 net6545 net6416 net6625 vdd vss unit_coupling_tile
xi1559 net6547 net6422 net6549 net6548 net6545 net6550 net6421 net6546 vdd vss unit_coupling_tile
xi1558 net6557 net6343 net6555 net6549 net6550 net6552 net6342 net6556 vdd vss unit_coupling_tile
xi1557 net6554 net6353 net6563 net6555 net6552 net6560 net6352 net6553 vdd vss unit_coupling_tile
xi1556 net6562 net6350 net6564 net6563 net6560 net6558 net6349 net6561 vdd vss unit_coupling_tile
xi1555 net6571 net6358 net6568 net6564 net6558 net6565 net6357 net6559 vdd vss unit_coupling_tile
xi1554 net6567 net6367 net6569 net6568 net6565 net6570 net6355 net6566 vdd vss unit_coupling_tile
xi1553 net6576 net6363 net6577 net6569 net6570 net6572 net6362 net6575 vdd vss unit_coupling_tile
xi1552 net6574 net6372 net6581 net6577 net6572 net6578 net6371 net6573 vdd vss unit_coupling_tile
xi1551 net6580 net6370 net6582 net6581 net6578 net6583 net6369 net6579 vdd vss unit_coupling_tile
xi1550 net6585 net6376 net6510 net6582 net6583 net6511 net6375 net6584 vdd vss unit_coupling_tile
xi1549 net6508 net6381 net6509 net72 net72 net6505 net6380 net6507 vdd vss unit_coupling_tile
xi1548 net6518 net6305 net6515 net6509 net6505 net6512 net6304 net6506 vdd vss unit_coupling_tile
xi1547 net6514 net6314 net6516 net6515 net6512 net6517 net6302 net6513 vdd vss unit_coupling_tile
xi1546 net6523 net6310 net6524 net6516 net6517 net6519 net6309 net6522 vdd vss unit_coupling_tile
xi1545 net6521 net6319 net6528 net6524 net6519 net6525 net6318 net6520 vdd vss unit_coupling_tile
xi1544 net6527 net6317 net6529 net6528 net6525 net6530 net6316 net6526 vdd vss unit_coupling_tile
xi1543 net6536 net6323 net6534 net6529 net6530 net6531 net6322 net6535 vdd vss unit_coupling_tile
xi1542 net6533 net6332 net6542 net6534 net6531 net6539 net6331 net6532 vdd vss unit_coupling_tile
xi1541 net6541 net6329 net6543 net6542 net6539 net6537 net6328 net6540 vdd vss unit_coupling_tile
xi1540 net6544 net6337 net6471 net6543 net6537 net6468 net6336 net6538 vdd vss unit_coupling_tile
xi1539 net6470 net6340 net6472 net6471 net6468 net6465 net6334 net6469 vdd vss unit_coupling_tile
xi1538 net6467 net6266 net6476 net6472 net6465 net6473 net6265 net6466 vdd vss unit_coupling_tile
xi1537 net6475 net6263 net6477 net6476 net6473 net6478 net6262 net6474 vdd vss unit_coupling_tile
xi1536 net6484 net6271 net6482 net6477 net6478 net6479 net6270 net6483 vdd vss unit_coupling_tile
xi1535 net6481 net6280 net6490 net6482 net6479 net6487 net6279 net6480 vdd vss unit_coupling_tile
xi1534 net6489 net6277 net6491 net6490 net6487 net6485 net6276 net6488 vdd vss unit_coupling_tile
xi1533 net6498 net6285 net6495 net6491 net6485 net6492 net6284 net6486 vdd vss unit_coupling_tile
xi1532 net6494 net6294 net6496 net6495 net6492 net6497 net6282 net6493 vdd vss unit_coupling_tile
xi1531 net6503 net6290 net6504 net6496 net6497 net6499 net6289 net6502 vdd vss unit_coupling_tile
xi1530 net6501 net6299 net6430 net6504 net6499 net6427 net6298 net6500 vdd vss unit_coupling_tile
xi1529 net6429 net6297 net6426 net6430 net6427 net6423 net6296 net6428 vdd vss unit_coupling_tile
xi1528 net6425 net6225 net6436 net6426 net6423 net6433 net6224 net6424 vdd vss unit_coupling_tile
xi1527 net6435 net6221 net6437 net6436 net6433 net6431 net6220 net6434 vdd vss unit_coupling_tile
xi1526 net6444 net6231 net6441 net6437 net6431 net6438 net6230 net6432 vdd vss unit_coupling_tile
xi1525 net6440 net6240 net6442 net6441 net6438 net6443 net6228 net6439 vdd vss unit_coupling_tile
xi1524 net6449 net6236 net6450 net6442 net6443 net6445 net6235 net6448 vdd vss unit_coupling_tile
xi1523 net6447 net6245 net6454 net6450 net6445 net6451 net6244 net6446 vdd vss unit_coupling_tile
xi1522 net6453 net6243 net6455 net6454 net6451 net6456 net6242 net6452 vdd vss unit_coupling_tile
xi1521 net6462 net6249 net6460 net6455 net6456 net6457 net6248 net6461 vdd vss unit_coupling_tile
xi1520 net6459 net6258 net6389 net6460 net6457 net6463 net6257 net6458 vdd vss unit_coupling_tile
xi1518 net6384 net6184 net6386 net6385 net6382 net6387 net6260 net6383 vdd vss unit_coupling_tile
xi1517 net6394 net6180 net6395 net6386 net6387 net6390 net6179 net6393 vdd vss unit_coupling_tile
xi1516 net6392 net6190 net6399 net6395 net6390 net6396 net6189 net6391 vdd vss unit_coupling_tile
xi1515 net6398 net6188 net6400 net6399 net6396 net6401 net6187 net6397 vdd vss unit_coupling_tile
xi1514 net6407 net6194 net6405 net6400 net6401 net6402 net6193 net6406 vdd vss unit_coupling_tile
xi1513 net6404 net6203 net6413 net6405 net6402 net6410 net6202 net6403 vdd vss unit_coupling_tile
xi1512 net6412 net6200 net6414 net6413 net6410 net6408 net6199 net6411 vdd vss unit_coupling_tile
xi1511 net6420 net6208 net6418 net6414 net6408 net6415 net6207 net6409 vdd vss unit_coupling_tile
xi1510 net6417 net6216 net6347 net6418 net6415 net6419 net6205 net6416 vdd vss unit_coupling_tile
xi1509 net6422 net6213 net6344 net6347 net6419 net6341 net6212 net6421 vdd vss unit_coupling_tile
xi1508 net6343 net6218 net6345 net6344 net6341 net6346 net6217 net6342 vdd vss unit_coupling_tile
xi1507 net6353 net6139 net6351 net6345 net6346 net6348 net6138 net6352 vdd vss unit_coupling_tile
xi1506 net6350 net6149 net6359 net6351 net6348 net6356 net6148 net6349 vdd vss unit_coupling_tile
xi1505 net6358 net6146 net6360 net6359 net6356 net6354 net6145 net6357 vdd vss unit_coupling_tile
xi1504 net6367 net6154 net6364 net6360 net6354 net6361 net6153 net6355 vdd vss unit_coupling_tile
xi1503 net6363 net6163 net6365 net6364 net6361 net6366 net6151 net6362 vdd vss unit_coupling_tile
xi1502 net6372 net6159 net6373 net6365 net6366 net6368 net6158 net6371 vdd vss unit_coupling_tile
xi1501 net6370 net6168 net6377 net6373 net6368 net6374 net6167 net6369 vdd vss unit_coupling_tile
xi1500 net6376 net6166 net6378 net6377 net6374 net6379 net6165 net6375 vdd vss unit_coupling_tile
xi1499 net6381 net6171 net6306 net73 net73 net6303 net6170 net6380 vdd vss unit_coupling_tile
xi1498 net6305 net6177 net6307 net6306 net6303 net6301 net6176 net6304 vdd vss unit_coupling_tile
xi1497 net6314 net6101 net6311 net6307 net6301 net6308 net6100 net6302 vdd vss unit_coupling_tile
xi1496 net6310 net6110 net6312 net6311 net6308 net6313 net6098 net6309 vdd vss unit_coupling_tile
xi1495 net6319 net6106 net6320 net6312 net6313 net6315 net6105 net6318 vdd vss unit_coupling_tile
xi1494 net6317 net6115 net6324 net6320 net6315 net6321 net6114 net6316 vdd vss unit_coupling_tile
xi1493 net6323 net6113 net6325 net6324 net6321 net6326 net6112 net6322 vdd vss unit_coupling_tile
xi1492 net6332 net6119 net6330 net6325 net6326 net6327 net6118 net6331 vdd vss unit_coupling_tile
xi1491 net6329 net6128 net6338 net6330 net6327 net6335 net6127 net6328 vdd vss unit_coupling_tile
xi1490 net6337 net6125 net6339 net6338 net6335 net6333 net6124 net6336 vdd vss unit_coupling_tile
xi1489 net6340 net6133 net6267 net6339 net6333 net6264 net6132 net6334 vdd vss unit_coupling_tile
xi1488 net6266 net6136 net6268 net6267 net6264 net6261 net6130 net6265 vdd vss unit_coupling_tile
xi1487 net6263 net6062 net6272 net6268 net6261 net6269 net6061 net6262 vdd vss unit_coupling_tile
xi1486 net6271 net6059 net6273 net6272 net6269 net6274 net6058 net6270 vdd vss unit_coupling_tile
xi1485 net6280 net6067 net6278 net6273 net6274 net6275 net6066 net6279 vdd vss unit_coupling_tile
xi1484 net6277 net6076 net6286 net6278 net6275 net6283 net6075 net6276 vdd vss unit_coupling_tile
xi1483 net6285 net6073 net6287 net6286 net6283 net6281 net6072 net6284 vdd vss unit_coupling_tile
xi1482 net6294 net6081 net6291 net6287 net6281 net6288 net6080 net6282 vdd vss unit_coupling_tile
xi1481 net6290 net6090 net6292 net6291 net6288 net6293 net6078 net6289 vdd vss unit_coupling_tile
xi1480 net6299 net6086 net6300 net6292 net6293 net6295 net6085 net6298 vdd vss unit_coupling_tile
xi1479 net6297 net6095 net6226 net6300 net6295 net6223 net6094 net6296 vdd vss unit_coupling_tile
xi1478 net6225 net6093 net6222 net6226 net6223 net6219 net6092 net6224 vdd vss unit_coupling_tile
xi1477 net6221 net6021 net6232 net6222 net6219 net6229 net6020 net6220 vdd vss unit_coupling_tile
xi1476 net6231 net6017 net6233 net6232 net6229 net6227 net6016 net6230 vdd vss unit_coupling_tile
xi1475 net6240 net6027 net6237 net6233 net6227 net6234 net6026 net6228 vdd vss unit_coupling_tile
xi1474 net6236 net6036 net6238 net6237 net6234 net6239 net6024 net6235 vdd vss unit_coupling_tile
xi1473 net6245 net6032 net6246 net6238 net6239 net6241 net6031 net6244 vdd vss unit_coupling_tile
xi1472 net6243 net6038 net6250 net6246 net6241 net6247 net6037 net6242 vdd vss unit_coupling_tile
xi1471 net6249 net6042 net6251 net6250 net6247 net6252 net6041 net6248 vdd vss unit_coupling_tile
xi1469 net6255 net6054 net6185 net6256 net6253 net6259 net6053 net6254 vdd vss unit_coupling_tile
xi1468 net6184 net6051 net6181 net6185 net6259 net6178 net6050 net6260 vdd vss unit_coupling_tile
xi1467 net6180 net5980 net6182 net6181 net6178 net6183 net6056 net6179 vdd vss unit_coupling_tile
xi1466 net6190 net5976 net6191 net6182 net6183 net6186 net5975 net6189 vdd vss unit_coupling_tile
xi1465 net6188 net5986 net6195 net6191 net6186 net6192 net5985 net6187 vdd vss unit_coupling_tile
xi1464 net6194 net5984 net6196 net6195 net6192 net6197 net5983 net6193 vdd vss unit_coupling_tile
xi1463 net6203 net5990 net6201 net6196 net6197 net6198 net5989 net6202 vdd vss unit_coupling_tile
xi1462 net6200 net5999 net6209 net6201 net6198 net6206 net5998 net6199 vdd vss unit_coupling_tile
xi1461 net6208 net5996 net6210 net6209 net6206 net6204 net5995 net6207 vdd vss unit_coupling_tile
xi1460 net6216 net6004 net6214 net6210 net6204 net6211 net6003 net6205 vdd vss unit_coupling_tile
xi1459 net6213 net6012 net6143 net6214 net6211 net6215 net6001 net6212 vdd vss unit_coupling_tile
xi1458 net6218 net6009 net6140 net6143 net6215 net6137 net6008 net6217 vdd vss unit_coupling_tile
xi1457 net6139 net6014 net6141 net6140 net6137 net6142 net6013 net6138 vdd vss unit_coupling_tile
xi1456 net6149 net5935 net6147 net6141 net6142 net6144 net5934 net6148 vdd vss unit_coupling_tile
xi1455 net6146 net5945 net6155 net6147 net6144 net6152 net5944 net6145 vdd vss unit_coupling_tile
xi1454 net6154 net5942 net6156 net6155 net6152 net6150 net5941 net6153 vdd vss unit_coupling_tile
xi1453 net6163 net5950 net6160 net6156 net6150 net6157 net5949 net6151 vdd vss unit_coupling_tile
xi1452 net6159 net5959 net6161 net6160 net6157 net6162 net5947 net6158 vdd vss unit_coupling_tile
xi1451 net6168 net5955 net6169 net6161 net6162 net6164 net5954 net6167 vdd vss unit_coupling_tile
xi1450 net6166 net5963 net6174 net6169 net6164 net6175 net5962 net6165 vdd vss unit_coupling_tile
xi1449 net6171 net5961 net6172 net74 net74 net6173 net5960 net6170 vdd vss unit_coupling_tile
xi1448 net6177 net5968 net6102 net6172 net6173 net6099 net5967 net6176 vdd vss unit_coupling_tile
xi1447 net6101 net5973 net6103 net6102 net6099 net6097 net5972 net6100 vdd vss unit_coupling_tile
xi1446 net6110 net5897 net6107 net6103 net6097 net6104 net5896 net6098 vdd vss unit_coupling_tile
xi1445 net6106 net5906 net6108 net6107 net6104 net6109 net5894 net6105 vdd vss unit_coupling_tile
xi1444 net6115 net5902 net6116 net6108 net6109 net6111 net5901 net6114 vdd vss unit_coupling_tile
xi1443 net6113 net5911 net6120 net6116 net6111 net6117 net5910 net6112 vdd vss unit_coupling_tile
xi1442 net6119 net5909 net6121 net6120 net6117 net6122 net5908 net6118 vdd vss unit_coupling_tile
xi1441 net6128 net5915 net6126 net6121 net6122 net6123 net5914 net6127 vdd vss unit_coupling_tile
xi1440 net6125 net5924 net6134 net6126 net6123 net6131 net5923 net6124 vdd vss unit_coupling_tile
xi1439 net6133 net5921 net6135 net6134 net6131 net6129 net5920 net6132 vdd vss unit_coupling_tile
xi1438 net6136 net5929 net6063 net6135 net6129 net6060 net5928 net6130 vdd vss unit_coupling_tile
xi1437 net6062 net5932 net6064 net6063 net6060 net6057 net5926 net6061 vdd vss unit_coupling_tile
xi1436 net6059 net5858 net6068 net6064 net6057 net6065 net5857 net6058 vdd vss unit_coupling_tile
xi1435 net6067 net5855 net6069 net6068 net6065 net6070 net5854 net6066 vdd vss unit_coupling_tile
xi1434 net6076 net5863 net6074 net6069 net6070 net6071 net5862 net6075 vdd vss unit_coupling_tile
xi1433 net6073 net5872 net6082 net6074 net6071 net6079 net5871 net6072 vdd vss unit_coupling_tile
xi1432 net6081 net5869 net6083 net6082 net6079 net6077 net5868 net6080 vdd vss unit_coupling_tile
xi1431 net6090 net5877 net6087 net6083 net6077 net6084 net5876 net6078 vdd vss unit_coupling_tile
xi1430 net6086 net5886 net6088 net6087 net6084 net6089 net5874 net6085 vdd vss unit_coupling_tile
xi1429 net6095 net5882 net6096 net6088 net6089 net6091 net5881 net6094 vdd vss unit_coupling_tile
xi1428 net6093 net5891 net6022 net6096 net6091 net6019 net5890 net6092 vdd vss unit_coupling_tile
xi1427 net6021 net5889 net6018 net6022 net6019 net6015 net5888 net6020 vdd vss unit_coupling_tile
xi1426 net6017 net5817 net6028 net6018 net6015 net6025 net5816 net6016 vdd vss unit_coupling_tile
xi1425 net6027 net5813 net6029 net6028 net6025 net6023 net5812 net6026 vdd vss unit_coupling_tile
xi1424 net6036 net5823 net6033 net6029 net6023 net6030 net5822 net6024 vdd vss unit_coupling_tile
xi1423 net6032 net5826 net6034 net6033 net6030 net6035 net5820 net6031 vdd vss unit_coupling_tile
xi1422 net6038 net5830 net6039 net6034 net6035 net6040 net5829 net6037 vdd vss unit_coupling_tile
xi1420 net6045 net5835 net6047 net6046 net6043 net6048 net5834 net6044 vdd vss unit_coupling_tile
xi1419 net6054 net5841 net6052 net6047 net6048 net6049 net5840 net6053 vdd vss unit_coupling_tile
xi1418 net6051 net5850 net5981 net6052 net6049 net6055 net5849 net6050 vdd vss unit_coupling_tile
xi1417 net5980 net5847 net5977 net5981 net6055 net5974 net5846 net6056 vdd vss unit_coupling_tile
xi1416 net5976 net5776 net5978 net5977 net5974 net5979 net5852 net5975 vdd vss unit_coupling_tile
xi1415 net5986 net5772 net5987 net5978 net5979 net5982 net5771 net5985 vdd vss unit_coupling_tile
xi1414 net5984 net5782 net5991 net5987 net5982 net5988 net5781 net5983 vdd vss unit_coupling_tile
xi1413 net5990 net5780 net5992 net5991 net5988 net5993 net5779 net5989 vdd vss unit_coupling_tile
xi1412 net5999 net5786 net5997 net5992 net5993 net5994 net5785 net5998 vdd vss unit_coupling_tile
xi1411 net5996 net5795 net6005 net5997 net5994 net6002 net5794 net5995 vdd vss unit_coupling_tile
xi1410 net6004 net5792 net6006 net6005 net6002 net6000 net5791 net6003 vdd vss unit_coupling_tile
xi1409 net6012 net5800 net6010 net6006 net6000 net6007 net5799 net6001 vdd vss unit_coupling_tile
xi1408 net6009 net5808 net5939 net6010 net6007 net6011 net5797 net6008 vdd vss unit_coupling_tile
xi1407 net6014 net5805 net5936 net5939 net6011 net5933 net5804 net6013 vdd vss unit_coupling_tile
xi1406 net5935 net5810 net5937 net5936 net5933 net5938 net5809 net5934 vdd vss unit_coupling_tile
xi1405 net5945 net5731 net5943 net5937 net5938 net5940 net5730 net5944 vdd vss unit_coupling_tile
xi1404 net5942 net5741 net5951 net5943 net5940 net5948 net5740 net5941 vdd vss unit_coupling_tile
xi1403 net5950 net5738 net5952 net5951 net5948 net5946 net5737 net5949 vdd vss unit_coupling_tile
xi1402 net5959 net5746 net5956 net5952 net5946 net5953 net5745 net5947 vdd vss unit_coupling_tile
xi1401 net5955 net5755 net5957 net5956 net5953 net5958 net5743 net5954 vdd vss unit_coupling_tile
xi1400 net5963 net5751 net5964 net5957 net5958 net5965 net5750 net5962 vdd vss unit_coupling_tile
xi1399 net5961 net5760 net5969 net75 net75 net5966 net5759 net5960 vdd vss unit_coupling_tile
xi1398 net5968 net5758 net5970 net5969 net5966 net5971 net5757 net5967 vdd vss unit_coupling_tile
xi1397 net5973 net5764 net5898 net5970 net5971 net5895 net5763 net5972 vdd vss unit_coupling_tile
xi1396 net5897 net5769 net5899 net5898 net5895 net5893 net5768 net5896 vdd vss unit_coupling_tile
xi1395 net5906 net5693 net5903 net5899 net5893 net5900 net5692 net5894 vdd vss unit_coupling_tile
xi1394 net5902 net5702 net5904 net5903 net5900 net5905 net5690 net5901 vdd vss unit_coupling_tile
xi1393 net5911 net5698 net5912 net5904 net5905 net5907 net5697 net5910 vdd vss unit_coupling_tile
xi1392 net5909 net5707 net5916 net5912 net5907 net5913 net5706 net5908 vdd vss unit_coupling_tile
xi1391 net5915 net5705 net5917 net5916 net5913 net5918 net5704 net5914 vdd vss unit_coupling_tile
xi1390 net5924 net5711 net5922 net5917 net5918 net5919 net5710 net5923 vdd vss unit_coupling_tile
xi1389 net5921 net5720 net5930 net5922 net5919 net5927 net5719 net5920 vdd vss unit_coupling_tile
xi1388 net5929 net5717 net5931 net5930 net5927 net5925 net5716 net5928 vdd vss unit_coupling_tile
xi1387 net5932 net5725 net5859 net5931 net5925 net5856 net5724 net5926 vdd vss unit_coupling_tile
xi1386 net5858 net5728 net5860 net5859 net5856 net5853 net5722 net5857 vdd vss unit_coupling_tile
xi1385 net5855 net5654 net5864 net5860 net5853 net5861 net5653 net5854 vdd vss unit_coupling_tile
xi1384 net5863 net5651 net5865 net5864 net5861 net5866 net5650 net5862 vdd vss unit_coupling_tile
xi1383 net5872 net5659 net5870 net5865 net5866 net5867 net5658 net5871 vdd vss unit_coupling_tile
xi1382 net5869 net5668 net5878 net5870 net5867 net5875 net5667 net5868 vdd vss unit_coupling_tile
xi1381 net5877 net5665 net5879 net5878 net5875 net5873 net5664 net5876 vdd vss unit_coupling_tile
xi1380 net5886 net5673 net5883 net5879 net5873 net5880 net5672 net5874 vdd vss unit_coupling_tile
xi1379 net5882 net5682 net5884 net5883 net5880 net5885 net5670 net5881 vdd vss unit_coupling_tile
xi1378 net5891 net5678 net5892 net5884 net5885 net5887 net5677 net5890 vdd vss unit_coupling_tile
xi1377 net5889 net5687 net5818 net5892 net5887 net5815 net5686 net5888 vdd vss unit_coupling_tile
xi1376 net5817 net5685 net5814 net5818 net5815 net5811 net5684 net5816 vdd vss unit_coupling_tile
xi1375 net5813 net5613 net5824 net5814 net5811 net5821 net5612 net5812 vdd vss unit_coupling_tile
xi1374 net5823 net5609 net5825 net5824 net5821 net5819 net5608 net5822 vdd vss unit_coupling_tile
xi1373 net5826 net5620 net5827 net5825 net5819 net5828 net5619 net5820 vdd vss unit_coupling_tile
xi1371 net5837 net5624 net5838 net5831 net5832 net5833 net5623 net5836 vdd vss unit_coupling_tile
xi1370 net5835 net5633 net5842 net5838 net5833 net5839 net5632 net5834 vdd vss unit_coupling_tile
xi1369 net5841 net5631 net5843 net5842 net5839 net5844 net5630 net5840 vdd vss unit_coupling_tile
xi1368 net5850 net5637 net5848 net5843 net5844 net5845 net5636 net5849 vdd vss unit_coupling_tile
xi1367 net5847 net5646 net5777 net5848 net5845 net5851 net5645 net5846 vdd vss unit_coupling_tile
xi1366 net5776 net5643 net5773 net5777 net5851 net5770 net5642 net5852 vdd vss unit_coupling_tile
xi1365 net5772 net5572 net5774 net5773 net5770 net5775 net5648 net5771 vdd vss unit_coupling_tile
xi1364 net5782 net5568 net5783 net5774 net5775 net5778 net5567 net5781 vdd vss unit_coupling_tile
xi1363 net5780 net5578 net5787 net5783 net5778 net5784 net5577 net5779 vdd vss unit_coupling_tile
xi1362 net5786 net5576 net5788 net5787 net5784 net5789 net5575 net5785 vdd vss unit_coupling_tile
xi1361 net5795 net5582 net5793 net5788 net5789 net5790 net5581 net5794 vdd vss unit_coupling_tile
xi1360 net5792 net5591 net5801 net5793 net5790 net5798 net5590 net5791 vdd vss unit_coupling_tile
xi1359 net5800 net5588 net5802 net5801 net5798 net5796 net5587 net5799 vdd vss unit_coupling_tile
xi1358 net5808 net5596 net5806 net5802 net5796 net5803 net5595 net5797 vdd vss unit_coupling_tile
xi1357 net5805 net5604 net5735 net5806 net5803 net5807 net5593 net5804 vdd vss unit_coupling_tile
xi1356 net5810 net5601 net5732 net5735 net5807 net5729 net5600 net5809 vdd vss unit_coupling_tile
xi1355 net5731 net5606 net5733 net5732 net5729 net5734 net5605 net5730 vdd vss unit_coupling_tile
xi1354 net5741 net5527 net5739 net5733 net5734 net5736 net5526 net5740 vdd vss unit_coupling_tile
xi1353 net5738 net5537 net5747 net5739 net5736 net5744 net5536 net5737 vdd vss unit_coupling_tile
xi1352 net5746 net5534 net5748 net5747 net5744 net5742 net5533 net5745 vdd vss unit_coupling_tile
xi1351 net5755 net5542 net5752 net5748 net5742 net5749 net5541 net5743 vdd vss unit_coupling_tile
xi1350 net5751 net5549 net5753 net5752 net5749 net5754 net5539 net5750 vdd vss unit_coupling_tile
xi1349 net5760 net5546 net5761 net76 net76 net5756 net5545 net5759 vdd vss unit_coupling_tile
xi1348 net5758 net5556 net5765 net5761 net5756 net5762 net5555 net5757 vdd vss unit_coupling_tile
xi1347 net5764 net5554 net5766 net5765 net5762 net5767 net5553 net5763 vdd vss unit_coupling_tile
xi1346 net5769 net5560 net5694 net5766 net5767 net5691 net5559 net5768 vdd vss unit_coupling_tile
xi1345 net5693 net5565 net5695 net5694 net5691 net5689 net5564 net5692 vdd vss unit_coupling_tile
xi1344 net5702 net5489 net5699 net5695 net5689 net5696 net5488 net5690 vdd vss unit_coupling_tile
xi1343 net5698 net5498 net5700 net5699 net5696 net5701 net5486 net5697 vdd vss unit_coupling_tile
xi1342 net5707 net5494 net5708 net5700 net5701 net5703 net5493 net5706 vdd vss unit_coupling_tile
xi1341 net5705 net5503 net5712 net5708 net5703 net5709 net5502 net5704 vdd vss unit_coupling_tile
xi1340 net5711 net5501 net5713 net5712 net5709 net5714 net5500 net5710 vdd vss unit_coupling_tile
xi1339 net5720 net5507 net5718 net5713 net5714 net5715 net5506 net5719 vdd vss unit_coupling_tile
xi1338 net5717 net5516 net5726 net5718 net5715 net5723 net5515 net5716 vdd vss unit_coupling_tile
xi1337 net5725 net5513 net5727 net5726 net5723 net5721 net5512 net5724 vdd vss unit_coupling_tile
xi1336 net5728 net5521 net5655 net5727 net5721 net5652 net5520 net5722 vdd vss unit_coupling_tile
xi1335 net5654 net5524 net5656 net5655 net5652 net5649 net5518 net5653 vdd vss unit_coupling_tile
xi1334 net5651 net5450 net5660 net5656 net5649 net5657 net5449 net5650 vdd vss unit_coupling_tile
xi1333 net5659 net5447 net5661 net5660 net5657 net5662 net5446 net5658 vdd vss unit_coupling_tile
xi1332 net5668 net5455 net5666 net5661 net5662 net5663 net5454 net5667 vdd vss unit_coupling_tile
xi1331 net5665 net5464 net5674 net5666 net5663 net5671 net5463 net5664 vdd vss unit_coupling_tile
xi1330 net5673 net5461 net5675 net5674 net5671 net5669 net5460 net5672 vdd vss unit_coupling_tile
xi1329 net5682 net5469 net5679 net5675 net5669 net5676 net5468 net5670 vdd vss unit_coupling_tile
xi1328 net5678 net5478 net5680 net5679 net5676 net5681 net5466 net5677 vdd vss unit_coupling_tile
xi1327 net5687 net5474 net5688 net5680 net5681 net5683 net5473 net5686 vdd vss unit_coupling_tile
xi1326 net5685 net5483 net5614 net5688 net5683 net5611 net5482 net5684 vdd vss unit_coupling_tile
xi1325 net5613 net5481 net5610 net5614 net5611 net5607 net5480 net5612 vdd vss unit_coupling_tile
xi1324 net5609 net5409 net5617 net5610 net5607 net5618 net5408 net5608 vdd vss unit_coupling_tile
xi1322 net5628 net5415 net5625 net5621 net5615 net5622 net5414 net5616 vdd vss unit_coupling_tile
xi1321 net5624 net5424 net5626 net5625 net5622 net5627 net5412 net5623 vdd vss unit_coupling_tile
xi1320 net5633 net5420 net5634 net5626 net5627 net5629 net5419 net5632 vdd vss unit_coupling_tile
xi1319 net5631 net5429 net5638 net5634 net5629 net5635 net5428 net5630 vdd vss unit_coupling_tile
xi1318 net5637 net5427 net5639 net5638 net5635 net5640 net5426 net5636 vdd vss unit_coupling_tile
xi1317 net5646 net5433 net5644 net5639 net5640 net5641 net5432 net5645 vdd vss unit_coupling_tile
xi1316 net5643 net5442 net5573 net5644 net5641 net5647 net5441 net5642 vdd vss unit_coupling_tile
xi1315 net5572 net5439 net5569 net5573 net5647 net5566 net5438 net5648 vdd vss unit_coupling_tile
xi1314 net5568 net5368 net5570 net5569 net5566 net5571 net5444 net5567 vdd vss unit_coupling_tile
xi1313 net5578 net5364 net5579 net5570 net5571 net5574 net5363 net5577 vdd vss unit_coupling_tile
xi1312 net5576 net5374 net5583 net5579 net5574 net5580 net5373 net5575 vdd vss unit_coupling_tile
xi1311 net5582 net5372 net5584 net5583 net5580 net5585 net5371 net5581 vdd vss unit_coupling_tile
xi1310 net5591 net5378 net5589 net5584 net5585 net5586 net5377 net5590 vdd vss unit_coupling_tile
xi1309 net5588 net5387 net5597 net5589 net5586 net5594 net5386 net5587 vdd vss unit_coupling_tile
xi1308 net5596 net5384 net5598 net5597 net5594 net5592 net5383 net5595 vdd vss unit_coupling_tile
xi1307 net5604 net5392 net5602 net5598 net5592 net5599 net5391 net5593 vdd vss unit_coupling_tile
xi1306 net5601 net5400 net5531 net5602 net5599 net5603 net5389 net5600 vdd vss unit_coupling_tile
xi1305 net5606 net5397 net5528 net5531 net5603 net5525 net5396 net5605 vdd vss unit_coupling_tile
xi1304 net5527 net5402 net5529 net5528 net5525 net5530 net5401 net5526 vdd vss unit_coupling_tile
xi1303 net5537 net5323 net5535 net5529 net5530 net5532 net5322 net5536 vdd vss unit_coupling_tile
xi1302 net5534 net5333 net5543 net5535 net5532 net5540 net5332 net5533 vdd vss unit_coupling_tile
xi1301 net5542 net5330 net5544 net5543 net5540 net5538 net5329 net5541 vdd vss unit_coupling_tile
xi1300 net5549 net5337 net5550 net5544 net5538 net5551 net5336 net5539 vdd vss unit_coupling_tile
xi1299 net5546 net5347 net5547 net77 net77 net5548 net5334 net5545 vdd vss unit_coupling_tile
xi1298 net5556 net5343 net5557 net5547 net5548 net5552 net5342 net5555 vdd vss unit_coupling_tile
xi1297 net5554 net5352 net5561 net5557 net5552 net5558 net5351 net5553 vdd vss unit_coupling_tile
xi1296 net5560 net5350 net5562 net5561 net5558 net5563 net5349 net5559 vdd vss unit_coupling_tile
xi1295 net5565 net5356 net5490 net5562 net5563 net5487 net5355 net5564 vdd vss unit_coupling_tile
xi1294 net5489 net5361 net5491 net5490 net5487 net5485 net5360 net5488 vdd vss unit_coupling_tile
xi1293 net5498 net5285 net5495 net5491 net5485 net5492 net5284 net5486 vdd vss unit_coupling_tile
xi1292 net5494 net5294 net5496 net5495 net5492 net5497 net5282 net5493 vdd vss unit_coupling_tile
xi1291 net5503 net5290 net5504 net5496 net5497 net5499 net5289 net5502 vdd vss unit_coupling_tile
xi1290 net5501 net5299 net5508 net5504 net5499 net5505 net5298 net5500 vdd vss unit_coupling_tile
xi1289 net5507 net5297 net5509 net5508 net5505 net5510 net5296 net5506 vdd vss unit_coupling_tile
xi1288 net5516 net5303 net5514 net5509 net5510 net5511 net5302 net5515 vdd vss unit_coupling_tile
xi1287 net5513 net5312 net5522 net5514 net5511 net5519 net5311 net5512 vdd vss unit_coupling_tile
xi1286 net5521 net5309 net5523 net5522 net5519 net5517 net5308 net5520 vdd vss unit_coupling_tile
xi1285 net5524 net5317 net5451 net5523 net5517 net5448 net5316 net5518 vdd vss unit_coupling_tile
xi1284 net5450 net5320 net5452 net5451 net5448 net5445 net5314 net5449 vdd vss unit_coupling_tile
xi1283 net5447 net5246 net5456 net5452 net5445 net5453 net5245 net5446 vdd vss unit_coupling_tile
xi1282 net5455 net5243 net5457 net5456 net5453 net5458 net5242 net5454 vdd vss unit_coupling_tile
xi1281 net5464 net5251 net5462 net5457 net5458 net5459 net5250 net5463 vdd vss unit_coupling_tile
xi1280 net5461 net5260 net5470 net5462 net5459 net5467 net5259 net5460 vdd vss unit_coupling_tile
xi1279 net5469 net5257 net5471 net5470 net5467 net5465 net5256 net5468 vdd vss unit_coupling_tile
xi1278 net5478 net5265 net5475 net5471 net5465 net5472 net5264 net5466 vdd vss unit_coupling_tile
xi1277 net5474 net5274 net5476 net5475 net5472 net5477 net5262 net5473 vdd vss unit_coupling_tile
xi1276 net5483 net5270 net5484 net5476 net5477 net5479 net5269 net5482 vdd vss unit_coupling_tile
xi1275 net5481 net5279 net5410 net5484 net5479 net5407 net5278 net5480 vdd vss unit_coupling_tile
xi1273 net5405 net5205 net5416 net5406 net5403 net5413 net5204 net5404 vdd vss unit_coupling_tile
xi1272 net5415 net5201 net5417 net5416 net5413 net5411 net5200 net5414 vdd vss unit_coupling_tile
xi1271 net5424 net5211 net5421 net5417 net5411 net5418 net5210 net5412 vdd vss unit_coupling_tile
xi1270 net5420 net5220 net5422 net5421 net5418 net5423 net5208 net5419 vdd vss unit_coupling_tile
xi1269 net5429 net5216 net5430 net5422 net5423 net5425 net5215 net5428 vdd vss unit_coupling_tile
xi1268 net5427 net5225 net5434 net5430 net5425 net5431 net5224 net5426 vdd vss unit_coupling_tile
xi1267 net5433 net5223 net5435 net5434 net5431 net5436 net5222 net5432 vdd vss unit_coupling_tile
xi1266 net5442 net5229 net5440 net5435 net5436 net5437 net5228 net5441 vdd vss unit_coupling_tile
xi1265 net5439 net5238 net5369 net5440 net5437 net5443 net5237 net5438 vdd vss unit_coupling_tile
xi1264 net5368 net5235 net5365 net5369 net5443 net5362 net5234 net5444 vdd vss unit_coupling_tile
xi1263 net5364 net5164 net5366 net5365 net5362 net5367 net5240 net5363 vdd vss unit_coupling_tile
xi1262 net5374 net5160 net5375 net5366 net5367 net5370 net5159 net5373 vdd vss unit_coupling_tile
xi1261 net5372 net5170 net5379 net5375 net5370 net5376 net5169 net5371 vdd vss unit_coupling_tile
xi1260 net5378 net5168 net5380 net5379 net5376 net5381 net5167 net5377 vdd vss unit_coupling_tile
xi1259 net5387 net5174 net5385 net5380 net5381 net5382 net5173 net5386 vdd vss unit_coupling_tile
xi1258 net5384 net5183 net5393 net5385 net5382 net5390 net5182 net5383 vdd vss unit_coupling_tile
xi1257 net5392 net5180 net5394 net5393 net5390 net5388 net5179 net5391 vdd vss unit_coupling_tile
xi1256 net5400 net5188 net5398 net5394 net5388 net5395 net5187 net5389 vdd vss unit_coupling_tile
xi1255 net5397 net5196 net5327 net5398 net5395 net5399 net5185 net5396 vdd vss unit_coupling_tile
xi1254 net5402 net5193 net5324 net5327 net5399 net5321 net5192 net5401 vdd vss unit_coupling_tile
xi1253 net5323 net5198 net5325 net5324 net5321 net5326 net5197 net5322 vdd vss unit_coupling_tile
xi1252 net5333 net5119 net5331 net5325 net5326 net5328 net5118 net5332 vdd vss unit_coupling_tile
xi1251 net5330 net5129 net5338 net5331 net5328 net5335 net5128 net5329 vdd vss unit_coupling_tile
xi1250 net5337 net5126 net5339 net5338 net5335 net5340 net5125 net5336 vdd vss unit_coupling_tile
xi1249 net5347 net5133 net5344 net78 net78 net5341 net5132 net5334 vdd vss unit_coupling_tile
xi1248 net5343 net5143 net5345 net5344 net5341 net5346 net5131 net5342 vdd vss unit_coupling_tile
xi1247 net5352 net5139 net5353 net5345 net5346 net5348 net5138 net5351 vdd vss unit_coupling_tile
xi1246 net5350 net5148 net5357 net5353 net5348 net5354 net5147 net5349 vdd vss unit_coupling_tile
xi1245 net5356 net5146 net5358 net5357 net5354 net5359 net5145 net5355 vdd vss unit_coupling_tile
xi1244 net5361 net5152 net5286 net5358 net5359 net5283 net5151 net5360 vdd vss unit_coupling_tile
xi1243 net5285 net5157 net5287 net5286 net5283 net5281 net5156 net5284 vdd vss unit_coupling_tile
xi1242 net5294 net5081 net5291 net5287 net5281 net5288 net5080 net5282 vdd vss unit_coupling_tile
xi1241 net5290 net5090 net5292 net5291 net5288 net5293 net5078 net5289 vdd vss unit_coupling_tile
xi1240 net5299 net5086 net5300 net5292 net5293 net5295 net5085 net5298 vdd vss unit_coupling_tile
xi1239 net5297 net5095 net5304 net5300 net5295 net5301 net5094 net5296 vdd vss unit_coupling_tile
xi1238 net5303 net5093 net5305 net5304 net5301 net5306 net5092 net5302 vdd vss unit_coupling_tile
xi1237 net5312 net5099 net5310 net5305 net5306 net5307 net5098 net5311 vdd vss unit_coupling_tile
xi1236 net5309 net5108 net5318 net5310 net5307 net5315 net5107 net5308 vdd vss unit_coupling_tile
xi1235 net5317 net5105 net5319 net5318 net5315 net5313 net5104 net5316 vdd vss unit_coupling_tile
xi1234 net5320 net5113 net5247 net5319 net5313 net5244 net5112 net5314 vdd vss unit_coupling_tile
xi1233 net5246 net5116 net5248 net5247 net5244 net5241 net5110 net5245 vdd vss unit_coupling_tile
xi1232 net5243 net5042 net5252 net5248 net5241 net5249 net5041 net5242 vdd vss unit_coupling_tile
xi1231 net5251 net5039 net5253 net5252 net5249 net5254 net5038 net5250 vdd vss unit_coupling_tile
xi1230 net5260 net5047 net5258 net5253 net5254 net5255 net5046 net5259 vdd vss unit_coupling_tile
xi1229 net5257 net5056 net5266 net5258 net5255 net5263 net5055 net5256 vdd vss unit_coupling_tile
xi1228 net5265 net5053 net5267 net5266 net5263 net5261 net5052 net5264 vdd vss unit_coupling_tile
xi1227 net5274 net5059 net5271 net5267 net5261 net5268 net5058 net5262 vdd vss unit_coupling_tile
xi1226 net5270 net5070 net5272 net5271 net5268 net5273 net5063 net5269 vdd vss unit_coupling_tile
xi1224 net5277 net5075 net5206 net5280 net5275 net5203 net5074 net5276 vdd vss unit_coupling_tile
xi1223 net5205 net5073 net5202 net5206 net5203 net5199 net5072 net5204 vdd vss unit_coupling_tile
xi1222 net5201 net5001 net5212 net5202 net5199 net5209 net5000 net5200 vdd vss unit_coupling_tile
xi1221 net5211 net4997 net5213 net5212 net5209 net5207 net4996 net5210 vdd vss unit_coupling_tile
xi1220 net5220 net5007 net5217 net5213 net5207 net5214 net5006 net5208 vdd vss unit_coupling_tile
xi1219 net5216 net5016 net5218 net5217 net5214 net5219 net5004 net5215 vdd vss unit_coupling_tile
xi1218 net5225 net5012 net5226 net5218 net5219 net5221 net5011 net5224 vdd vss unit_coupling_tile
xi1217 net5223 net5021 net5230 net5226 net5221 net5227 net5020 net5222 vdd vss unit_coupling_tile
xi1216 net5229 net5019 net5231 net5230 net5227 net5232 net5018 net5228 vdd vss unit_coupling_tile
xi1215 net5238 net5025 net5236 net5231 net5232 net5233 net5024 net5237 vdd vss unit_coupling_tile
xi1214 net5235 net5034 net5165 net5236 net5233 net5239 net5033 net5234 vdd vss unit_coupling_tile
xi1213 net5164 net5031 net5161 net5165 net5239 net5158 net5030 net5240 vdd vss unit_coupling_tile
xi1212 net5160 net4960 net5162 net5161 net5158 net5163 net5036 net5159 vdd vss unit_coupling_tile
xi1211 net5170 net4956 net5171 net5162 net5163 net5166 net4955 net5169 vdd vss unit_coupling_tile
xi1210 net5168 net4966 net5175 net5171 net5166 net5172 net4965 net5167 vdd vss unit_coupling_tile
xi1209 net5174 net4964 net5176 net5175 net5172 net5177 net4963 net5173 vdd vss unit_coupling_tile
xi1208 net5183 net4970 net5181 net5176 net5177 net5178 net4969 net5182 vdd vss unit_coupling_tile
xi1207 net5180 net4979 net5189 net5181 net5178 net5186 net4978 net5179 vdd vss unit_coupling_tile
xi1206 net5188 net4976 net5190 net5189 net5186 net5184 net4975 net5187 vdd vss unit_coupling_tile
xi1205 net5196 net4984 net5194 net5190 net5184 net5191 net4983 net5185 vdd vss unit_coupling_tile
xi1204 net5193 net4992 net5123 net5194 net5191 net5195 net4981 net5192 vdd vss unit_coupling_tile
xi1203 net5198 net4989 net5120 net5123 net5195 net5117 net4988 net5197 vdd vss unit_coupling_tile
xi1202 net5119 net4994 net5121 net5120 net5117 net5122 net4993 net5118 vdd vss unit_coupling_tile
xi1201 net5129 net4915 net5127 net5121 net5122 net5124 net4914 net5128 vdd vss unit_coupling_tile
xi1200 net5126 net4923 net5135 net5127 net5124 net5136 net4922 net5125 vdd vss unit_coupling_tile
xi1199 net5133 net4921 net5134 net79 net79 net5130 net4920 net5132 vdd vss unit_coupling_tile
xi1198 net5143 net4930 net5140 net5134 net5130 net5137 net4929 net5131 vdd vss unit_coupling_tile
xi1197 net5139 net4939 net5141 net5140 net5137 net5142 net4927 net5138 vdd vss unit_coupling_tile
xi1196 net5148 net4935 net5149 net5141 net5142 net5144 net4934 net5147 vdd vss unit_coupling_tile
xi1195 net5146 net4944 net5153 net5149 net5144 net5150 net4943 net5145 vdd vss unit_coupling_tile
xi1194 net5152 net4942 net5154 net5153 net5150 net5155 net4941 net5151 vdd vss unit_coupling_tile
xi1193 net5157 net4948 net5082 net5154 net5155 net5079 net4947 net5156 vdd vss unit_coupling_tile
xi1192 net5081 net4953 net5083 net5082 net5079 net5077 net4952 net5080 vdd vss unit_coupling_tile
xi1191 net5090 net4877 net5087 net5083 net5077 net5084 net4876 net5078 vdd vss unit_coupling_tile
xi1190 net5086 net4886 net5088 net5087 net5084 net5089 net4874 net5085 vdd vss unit_coupling_tile
xi1189 net5095 net4882 net5096 net5088 net5089 net5091 net4881 net5094 vdd vss unit_coupling_tile
xi1188 net5093 net4891 net5100 net5096 net5091 net5097 net4890 net5092 vdd vss unit_coupling_tile
xi1187 net5099 net4889 net5101 net5100 net5097 net5102 net4888 net5098 vdd vss unit_coupling_tile
xi1186 net5108 net4895 net5106 net5101 net5102 net5103 net4894 net5107 vdd vss unit_coupling_tile
xi1185 net5105 net4904 net5114 net5106 net5103 net5111 net4903 net5104 vdd vss unit_coupling_tile
xi1184 net5113 net4901 net5115 net5114 net5111 net5109 net4900 net5112 vdd vss unit_coupling_tile
xi1183 net5116 net4909 net5043 net5115 net5109 net5040 net4908 net5110 vdd vss unit_coupling_tile
xi1182 net5042 net4912 net5044 net5043 net5040 net5037 net4906 net5041 vdd vss unit_coupling_tile
xi1181 net5039 net4838 net5048 net5044 net5037 net5045 net4837 net5038 vdd vss unit_coupling_tile
xi1180 net5047 net4835 net5049 net5048 net5045 net5050 net4834 net5046 vdd vss unit_coupling_tile
xi1179 net5056 net4843 net5054 net5049 net5050 net5051 net4842 net5055 vdd vss unit_coupling_tile
xi1178 net5053 net4848 net5060 net5054 net5051 net5057 net4847 net5052 vdd vss unit_coupling_tile
xi1177 net5059 net4852 net5061 net5060 net5057 net5062 net4851 net5058 vdd vss unit_coupling_tile
xi1175 net5066 net4866 net5068 net5067 net5064 net5069 net4854 net5065 vdd vss unit_coupling_tile
xi1174 net5075 net4862 net5076 net5068 net5069 net5071 net4861 net5074 vdd vss unit_coupling_tile
xi1173 net5073 net4871 net5002 net5076 net5071 net4999 net4870 net5072 vdd vss unit_coupling_tile
xi1172 net5001 net4869 net4998 net5002 net4999 net4995 net4868 net5000 vdd vss unit_coupling_tile
xi1171 net4997 net4797 net5008 net4998 net4995 net5005 net4796 net4996 vdd vss unit_coupling_tile
xi1170 net5007 net4793 net5009 net5008 net5005 net5003 net4792 net5006 vdd vss unit_coupling_tile
xi1169 net5016 net4803 net5013 net5009 net5003 net5010 net4802 net5004 vdd vss unit_coupling_tile
xi1168 net5012 net4812 net5014 net5013 net5010 net5015 net4800 net5011 vdd vss unit_coupling_tile
xi1167 net5021 net4808 net5022 net5014 net5015 net5017 net4807 net5020 vdd vss unit_coupling_tile
xi1166 net5019 net4815 net5026 net5022 net5017 net5023 net4816 net5018 vdd vss unit_coupling_tile
xi1165 net5025 net4817 net5027 net5026 net5023 net5028 net4818 net5024 vdd vss unit_coupling_tile
xi1164 net5034 net4823 net5032 net5027 net5028 net5029 net4824 net5033 vdd vss unit_coupling_tile
xi1163 net5031 net4827 net4961 net5032 net5029 net5035 net4828 net5030 vdd vss unit_coupling_tile
xi1162 net4960 net4829 net4957 net4961 net5035 net4954 net4830 net5036 vdd vss unit_coupling_tile
xi1161 net4956 net4753 net4958 net4957 net4954 net4959 net4832 net4955 vdd vss unit_coupling_tile
xi1160 net4966 net4756 net4967 net4958 net4959 net4962 net4757 net4965 vdd vss unit_coupling_tile
xi1159 net4964 net4760 net4971 net4967 net4962 net4968 net4761 net4963 vdd vss unit_coupling_tile
xi1158 net4970 net4762 net4972 net4971 net4968 net4973 net4763 net4969 vdd vss unit_coupling_tile
xi1157 net4979 net4768 net4977 net4972 net4973 net4974 net4769 net4978 vdd vss unit_coupling_tile
xi1156 net4976 net4772 net4985 net4977 net4974 net4982 net4773 net4975 vdd vss unit_coupling_tile
xi1155 net4984 net4774 net4986 net4985 net4982 net4980 net4775 net4983 vdd vss unit_coupling_tile
xi1154 net4992 net4780 net4990 net4986 net4980 net4987 net4781 net4981 vdd vss unit_coupling_tile
xi1153 net4989 net4785 net4919 net4990 net4987 net4991 net4782 net4988 vdd vss unit_coupling_tile
xi1152 net4994 net4787 net4916 net4919 net4991 net4913 net4788 net4993 vdd vss unit_coupling_tile
xi1151 net4915 net4789 net4917 net4916 net4913 net4918 net4790 net4914 vdd vss unit_coupling_tile
xi1150 net4923 net4714 net4924 net4917 net4918 net4925 net4715 net4922 vdd vss unit_coupling_tile
xi1149 net4921 net4718 net4931 net80 net80 net4928 net4719 net4920 vdd vss unit_coupling_tile
xi1148 net4930 net4720 net4932 net4931 net4928 net4926 net4721 net4929 vdd vss unit_coupling_tile
xi1147 net4939 net4726 net4936 net4932 net4926 net4933 net4727 net4927 vdd vss unit_coupling_tile
xi1146 net4935 net4731 net4937 net4936 net4933 net4938 net4728 net4934 vdd vss unit_coupling_tile
xi1145 net4944 net4734 net4945 net4937 net4938 net4940 net4735 net4943 vdd vss unit_coupling_tile
xi1144 net4942 net4738 net4949 net4945 net4940 net4946 net4739 net4941 vdd vss unit_coupling_tile
xi1143 net4948 net4740 net4950 net4949 net4946 net4951 net4741 net4947 vdd vss unit_coupling_tile
xi1142 net4953 net4746 net4878 net4950 net4951 net4875 net4747 net4952 vdd vss unit_coupling_tile
xi1141 net4877 net4748 net4879 net4878 net4875 net4873 net4749 net4876 vdd vss unit_coupling_tile
xi1140 net4886 net4673 net4883 net4879 net4873 net4880 net4674 net4874 vdd vss unit_coupling_tile
xi1139 net4882 net4678 net4884 net4883 net4880 net4885 net4675 net4881 vdd vss unit_coupling_tile
xi1138 net4891 net4681 net4892 net4884 net4885 net4887 net4682 net4890 vdd vss unit_coupling_tile
xi1137 net4889 net4685 net4896 net4892 net4887 net4893 net4686 net4888 vdd vss unit_coupling_tile
xi1136 net4895 net4687 net4897 net4896 net4893 net4898 net4688 net4894 vdd vss unit_coupling_tile
xi1135 net4904 net4693 net4902 net4897 net4898 net4899 net4694 net4903 vdd vss unit_coupling_tile
xi1134 net4901 net4697 net4910 net4902 net4899 net4907 net4698 net4900 vdd vss unit_coupling_tile
xi1133 net4909 net4699 net4911 net4910 net4907 net4905 net4700 net4908 vdd vss unit_coupling_tile
xi1132 net4912 net4705 net4839 net4911 net4905 net4836 net4706 net4906 vdd vss unit_coupling_tile
xi1131 net4838 net4708 net4840 net4839 net4836 net4833 net4707 net4837 vdd vss unit_coupling_tile
xi1130 net4835 net4632 net4844 net4840 net4833 net4841 net4633 net4834 vdd vss unit_coupling_tile
xi1129 net4843 net4635 net4845 net4844 net4841 net4846 net4636 net4842 vdd vss unit_coupling_tile
xi1128 net4848 net4640 net4849 net4845 net4846 net4850 net4639 net4847 vdd vss unit_coupling_tile
xi1126 net4857 net4647 net4859 net4858 net4855 net4853 net4648 net4856 vdd vss unit_coupling_tile
xi1125 net4866 net4653 net4863 net4859 net4853 net4860 net4654 net4854 vdd vss unit_coupling_tile
xi1124 net4862 net4658 net4864 net4863 net4860 net4865 net4655 net4861 vdd vss unit_coupling_tile
xi1123 net4871 net4661 net4872 net4864 net4865 net4867 net4662 net4870 vdd vss unit_coupling_tile
xi1122 net4869 net4665 net4798 net4872 net4867 net4795 net4666 net4868 vdd vss unit_coupling_tile
xi1121 net4797 net4667 net4794 net4798 net4795 net4791 net4668 net4796 vdd vss unit_coupling_tile
xi1120 net4793 net4590 net4804 net4794 net4791 net4801 net4591 net4792 vdd vss unit_coupling_tile
xi1119 net4803 net4593 net4805 net4804 net4801 net4799 net4594 net4802 vdd vss unit_coupling_tile
xi1118 net4812 net4599 net4809 net4805 net4799 net4806 net4600 net4800 vdd vss unit_coupling_tile
xi1117 net4808 net4604 net4810 net4809 net4806 net4811 net4601 net4807 vdd vss unit_coupling_tile
xi1116 net4815 net4607 net4814 net4810 net4811 net4813 net4608 net4816 vdd vss unit_coupling_tile
xi1115 net4817 net4611 net4820 net4814 net4813 net4819 net4612 net4818 vdd vss unit_coupling_tile
xi1114 net4823 net4613 net4822 net4820 net4819 net4821 net4614 net4824 vdd vss unit_coupling_tile
xi1113 net4827 net4619 net4826 net4822 net4821 net4825 net4620 net4828 vdd vss unit_coupling_tile
xi1112 net4829 net4623 net4752 net4826 net4825 net4831 net4624 net4830 vdd vss unit_coupling_tile
xi1111 net4753 net4625 net4751 net4752 net4831 net4750 net4626 net4832 vdd vss unit_coupling_tile
xi1110 net4756 net4549 net4755 net4751 net4750 net4754 net4628 net4757 vdd vss unit_coupling_tile
xi1109 net4760 net4552 net4759 net4755 net4754 net4758 net4553 net4761 vdd vss unit_coupling_tile
xi1108 net4762 net4556 net4765 net4759 net4758 net4764 net4557 net4763 vdd vss unit_coupling_tile
xi1107 net4768 net4558 net4767 net4765 net4764 net4766 net4559 net4769 vdd vss unit_coupling_tile
xi1106 net4772 net4564 net4771 net4767 net4766 net4770 net4565 net4773 vdd vss unit_coupling_tile
xi1105 net4774 net4568 net4777 net4771 net4770 net4776 net4569 net4775 vdd vss unit_coupling_tile
xi1104 net4780 net4570 net4779 net4777 net4776 net4778 net4571 net4781 vdd vss unit_coupling_tile
xi1103 net4785 net4576 net4784 net4779 net4778 net4783 net4577 net4782 vdd vss unit_coupling_tile
xi1102 net4787 net4581 net4711 net4784 net4783 net4786 net4578 net4788 vdd vss unit_coupling_tile
xi1101 net4789 net4583 net4710 net4711 net4786 net4709 net4584 net4790 vdd vss unit_coupling_tile
xi1100 net4714 net4585 net4713 net4710 net4709 net4712 net4586 net4715 vdd vss unit_coupling_tile
xi1099 net4718 net4510 net4717 net81 net81 net4716 net4511 net4719 vdd vss unit_coupling_tile
xi1098 net4720 net4514 net4723 net4717 net4716 net4722 net4515 net4721 vdd vss unit_coupling_tile
xi1097 net4726 net4516 net4725 net4723 net4722 net4724 net4517 net4727 vdd vss unit_coupling_tile
xi1096 net4731 net4522 net4730 net4725 net4724 net4729 net4523 net4728 vdd vss unit_coupling_tile
xi1095 net4734 net4527 net4733 net4730 net4729 net4732 net4524 net4735 vdd vss unit_coupling_tile
xi1094 net4738 net4530 net4737 net4733 net4732 net4736 net4531 net4739 vdd vss unit_coupling_tile
xi1093 net4740 net4534 net4743 net4737 net4736 net4742 net4535 net4741 vdd vss unit_coupling_tile
xi1092 net4746 net4536 net4745 net4743 net4742 net4744 net4537 net4747 vdd vss unit_coupling_tile
xi1091 net4748 net4542 net4670 net4745 net4744 net4669 net4543 net4749 vdd vss unit_coupling_tile
xi1090 net4673 net4544 net4672 net4670 net4669 net4671 net4545 net4674 vdd vss unit_coupling_tile
xi1089 net4678 net4469 net4677 net4672 net4671 net4676 net4470 net4675 vdd vss unit_coupling_tile
xi1088 net4681 net4474 net4680 net4677 net4676 net4679 net4471 net4682 vdd vss unit_coupling_tile
xi1087 net4685 net4477 net4684 net4680 net4679 net4683 net4478 net4686 vdd vss unit_coupling_tile
xi1086 net4687 net4481 net4690 net4684 net4683 net4689 net4482 net4688 vdd vss unit_coupling_tile
xi1085 net4693 net4483 net4692 net4690 net4689 net4691 net4484 net4694 vdd vss unit_coupling_tile
xi1084 net4697 net4489 net4696 net4692 net4691 net4695 net4490 net4698 vdd vss unit_coupling_tile
xi1083 net4699 net4493 net4702 net4696 net4695 net4701 net4494 net4700 vdd vss unit_coupling_tile
xi1082 net4705 net4495 net4704 net4702 net4701 net4703 net4496 net4706 vdd vss unit_coupling_tile
xi1081 net4708 net4501 net4631 net4704 net4703 net4634 net4502 net4707 vdd vss unit_coupling_tile
xi1080 net4632 net4504 net4630 net4631 net4634 net4629 net4503 net4633 vdd vss unit_coupling_tile
xi1079 net4635 net4430 net4638 net4630 net4629 net4637 net4429 net4636 vdd vss unit_coupling_tile
xi1077 net4645 net4437 net4644 net4641 net4642 net4643 net4438 net4646 vdd vss unit_coupling_tile
xi1076 net4647 net4441 net4650 net4644 net4643 net4649 net4442 net4648 vdd vss unit_coupling_tile
xi1075 net4653 net4443 net4652 net4650 net4649 net4651 net4444 net4654 vdd vss unit_coupling_tile
xi1074 net4658 net4449 net4657 net4652 net4651 net4656 net4450 net4655 vdd vss unit_coupling_tile
xi1073 net4661 net4454 net4660 net4657 net4656 net4659 net4451 net4662 vdd vss unit_coupling_tile
xi1072 net4665 net4457 net4664 net4660 net4659 net4663 net4458 net4666 vdd vss unit_coupling_tile
xi1071 net4667 net4461 net4589 net4664 net4663 net4592 net4462 net4668 vdd vss unit_coupling_tile
xi1070 net4590 net4463 net4588 net4589 net4592 net4587 net4464 net4591 vdd vss unit_coupling_tile
xi1069 net4593 net4386 net4596 net4588 net4587 net4595 net4387 net4594 vdd vss unit_coupling_tile
xi1068 net4599 net4389 net4598 net4596 net4595 net4597 net4390 net4600 vdd vss unit_coupling_tile
xi1067 net4604 net4395 net4603 net4598 net4597 net4602 net4396 net4601 vdd vss unit_coupling_tile
xi1066 net4607 net4400 net4606 net4603 net4602 net4605 net4397 net4608 vdd vss unit_coupling_tile
xi1065 net4611 net4403 net4610 net4606 net4605 net4609 net4404 net4612 vdd vss unit_coupling_tile
xi1064 net4613 net4407 net4616 net4610 net4609 net4615 net4408 net4614 vdd vss unit_coupling_tile
xi1063 net4619 net4409 net4618 net4616 net4615 net4617 net4410 net4620 vdd vss unit_coupling_tile
xi1062 net4623 net4415 net4622 net4618 net4617 net4621 net4416 net4624 vdd vss unit_coupling_tile
xi1061 net4625 net4419 net4548 net4622 net4621 net4627 net4420 net4626 vdd vss unit_coupling_tile
xi1060 net4549 net4421 net4547 net4548 net4627 net4546 net4422 net4628 vdd vss unit_coupling_tile
xi1059 net4552 net4344 net4551 net4547 net4546 net4550 net4424 net4553 vdd vss unit_coupling_tile
xi1058 net4556 net4347 net4555 net4551 net4550 net4554 net4348 net4557 vdd vss unit_coupling_tile
xi1057 net4558 net4351 net4561 net4555 net4554 net4560 net4352 net4559 vdd vss unit_coupling_tile
xi1056 net4564 net4353 net4563 net4561 net4560 net4562 net4354 net4565 vdd vss unit_coupling_tile
xi1055 net4568 net4359 net4567 net4563 net4562 net4566 net4360 net4569 vdd vss unit_coupling_tile
xi1054 net4570 net4363 net4573 net4567 net4566 net4572 net4364 net4571 vdd vss unit_coupling_tile
xi1053 net4576 net4365 net4575 net4573 net4572 net4574 net4366 net4577 vdd vss unit_coupling_tile
xi1052 net4581 net4371 net4580 net4575 net4574 net4579 net4372 net4578 vdd vss unit_coupling_tile
xi1051 net4583 net4376 net4507 net4580 net4579 net4582 net4373 net4584 vdd vss unit_coupling_tile
xi1050 net4585 net4379 net4506 net4507 net4582 net4505 net4380 net4586 vdd vss unit_coupling_tile
xi1049 net4510 net4381 net4509 net82 net82 net4508 net4382 net4511 vdd vss unit_coupling_tile
xi1048 net4514 net4305 net4513 net4509 net4508 net4512 net4306 net4515 vdd vss unit_coupling_tile
xi1047 net4516 net4309 net4519 net4513 net4512 net4518 net4310 net4517 vdd vss unit_coupling_tile
xi1046 net4522 net4311 net4521 net4519 net4518 net4520 net4312 net4523 vdd vss unit_coupling_tile
xi1045 net4527 net4317 net4526 net4521 net4520 net4525 net4318 net4524 vdd vss unit_coupling_tile
xi1044 net4530 net4322 net4529 net4526 net4525 net4528 net4319 net4531 vdd vss unit_coupling_tile
xi1043 net4534 net4325 net4533 net4529 net4528 net4532 net4326 net4535 vdd vss unit_coupling_tile
xi1042 net4536 net4329 net4539 net4533 net4532 net4538 net4330 net4537 vdd vss unit_coupling_tile
xi1041 net4542 net4331 net4541 net4539 net4538 net4540 net4332 net4543 vdd vss unit_coupling_tile
xi1040 net4544 net4337 net4466 net4541 net4540 net4465 net4338 net4545 vdd vss unit_coupling_tile
xi1039 net4469 net4339 net4468 net4466 net4465 net4467 net4340 net4470 vdd vss unit_coupling_tile
xi1038 net4474 net4265 net4473 net4468 net4467 net4472 net4266 net4471 vdd vss unit_coupling_tile
xi1037 net4477 net4270 net4476 net4473 net4472 net4475 net4267 net4478 vdd vss unit_coupling_tile
xi1036 net4481 net4273 net4480 net4476 net4475 net4479 net4274 net4482 vdd vss unit_coupling_tile
xi1035 net4483 net4277 net4486 net4480 net4479 net4485 net4278 net4484 vdd vss unit_coupling_tile
xi1034 net4489 net4279 net4488 net4486 net4485 net4487 net4280 net4490 vdd vss unit_coupling_tile
xi1033 net4493 net4285 net4492 net4488 net4487 net4491 net4286 net4494 vdd vss unit_coupling_tile
xi1032 net4495 net4289 net4498 net4492 net4491 net4497 net4290 net4496 vdd vss unit_coupling_tile
xi1031 net4501 net4291 net4500 net4498 net4497 net4499 net4292 net4502 vdd vss unit_coupling_tile
xi1030 net4504 net4298 net4431 net4500 net4499 net4428 net4297 net4503 vdd vss unit_coupling_tile
xi1028 net4425 net4224 net4434 net4432 net4427 net4433 net4225 net4426 vdd vss unit_coupling_tile
xi1027 net4437 net4227 net4436 net4434 net4433 net4435 net4228 net4438 vdd vss unit_coupling_tile
xi1026 net4441 net4233 net4440 net4436 net4435 net4439 net4234 net4442 vdd vss unit_coupling_tile
xi1025 net4443 net4237 net4446 net4440 net4439 net4445 net4238 net4444 vdd vss unit_coupling_tile
xi1024 net4449 net4239 net4448 net4446 net4445 net4447 net4240 net4450 vdd vss unit_coupling_tile
xi1023 net4454 net4245 net4453 net4448 net4447 net4452 net4246 net4451 vdd vss unit_coupling_tile
xi1022 net4457 net4250 net4456 net4453 net4452 net4455 net4247 net4458 vdd vss unit_coupling_tile
xi1021 net4461 net4253 net4460 net4456 net4455 net4459 net4254 net4462 vdd vss unit_coupling_tile
xi1020 net4463 net4257 net4385 net4460 net4459 net4388 net4258 net4464 vdd vss unit_coupling_tile
xi1019 net4386 net4259 net4384 net4385 net4388 net4383 net4260 net4387 vdd vss unit_coupling_tile
xi1018 net4389 net4182 net4392 net4384 net4383 net4391 net4183 net4390 vdd vss unit_coupling_tile
xi1017 net4395 net4185 net4394 net4392 net4391 net4393 net4186 net4396 vdd vss unit_coupling_tile
xi1016 net4400 net4191 net4399 net4394 net4393 net4398 net4192 net4397 vdd vss unit_coupling_tile
xi1015 net4403 net4196 net4402 net4399 net4398 net4401 net4193 net4404 vdd vss unit_coupling_tile
xi1014 net4407 net4199 net4406 net4402 net4401 net4405 net4200 net4408 vdd vss unit_coupling_tile
xi1013 net4409 net4203 net4412 net4406 net4405 net4411 net4204 net4410 vdd vss unit_coupling_tile
xi1012 net4415 net4205 net4414 net4412 net4411 net4413 net4206 net4416 vdd vss unit_coupling_tile
xi1011 net4419 net4211 net4418 net4414 net4413 net4417 net4212 net4420 vdd vss unit_coupling_tile
xi1010 net4421 net4215 net4343 net4418 net4417 net4423 net4216 net4422 vdd vss unit_coupling_tile
xi1009 net4344 net4217 net4342 net4343 net4423 net4341 net4218 net4424 vdd vss unit_coupling_tile
xi1008 net4347 net4141 net4346 net4342 net4341 net4345 net4220 net4348 vdd vss unit_coupling_tile
xi1007 net4351 net4144 net4350 net4346 net4345 net4349 net4145 net4352 vdd vss unit_coupling_tile
xi1006 net4353 net4148 net4356 net4350 net4349 net4355 net4149 net4354 vdd vss unit_coupling_tile
xi1005 net4359 net4150 net4358 net4356 net4355 net4357 net4151 net4360 vdd vss unit_coupling_tile
xi1004 net4363 net4156 net4362 net4358 net4357 net4361 net4157 net4364 vdd vss unit_coupling_tile
xi1003 net4365 net4160 net4368 net4362 net4361 net4367 net4161 net4366 vdd vss unit_coupling_tile
xi1002 net4371 net4162 net4370 net4368 net4367 net4369 net4163 net4372 vdd vss unit_coupling_tile
xi1001 net4376 net4168 net4375 net4370 net4369 net4374 net4169 net4373 vdd vss unit_coupling_tile
xi1000 net4379 net4173 net4378 net4375 net4374 net4377 net4170 net4380 vdd vss unit_coupling_tile
xi999 net4381 net4175 net4302 net83 net83 net4301 net4176 net4382 vdd vss unit_coupling_tile
xi998 net4305 net4177 net4304 net4302 net4301 net4303 net4178 net4306 vdd vss unit_coupling_tile
xi997 net4309 net4102 net4308 net4304 net4303 net4307 net4103 net4310 vdd vss unit_coupling_tile
xi996 net4311 net4106 net4314 net4308 net4307 net4313 net4107 net4312 vdd vss unit_coupling_tile
xi995 net4317 net4108 net4316 net4314 net4313 net4315 net4109 net4318 vdd vss unit_coupling_tile
xi994 net4322 net4114 net4321 net4316 net4315 net4320 net4115 net4319 vdd vss unit_coupling_tile
xi993 net4325 net4119 net4324 net4321 net4320 net4323 net4116 net4326 vdd vss unit_coupling_tile
xi992 net4329 net4122 net4328 net4324 net4323 net4327 net4123 net4330 vdd vss unit_coupling_tile
xi991 net4331 net4126 net4334 net4328 net4327 net4333 net4127 net4332 vdd vss unit_coupling_tile
xi990 net4337 net4128 net4336 net4334 net4333 net4335 net4129 net4338 vdd vss unit_coupling_tile
xi989 net4339 net4134 net4262 net4336 net4335 net4261 net4135 net4340 vdd vss unit_coupling_tile
xi988 net4265 net4136 net4264 net4262 net4261 net4263 net4137 net4266 vdd vss unit_coupling_tile
xi987 net4270 net4061 net4269 net4264 net4263 net4268 net4062 net4267 vdd vss unit_coupling_tile
xi986 net4273 net4066 net4272 net4269 net4268 net4271 net4063 net4274 vdd vss unit_coupling_tile
xi985 net4277 net4069 net4276 net4272 net4271 net4275 net4070 net4278 vdd vss unit_coupling_tile
xi984 net4279 net4073 net4282 net4276 net4275 net4281 net4074 net4280 vdd vss unit_coupling_tile
xi983 net4285 net4075 net4284 net4282 net4281 net4283 net4076 net4286 vdd vss unit_coupling_tile
xi982 net4289 net4081 net4288 net4284 net4283 net4287 net4082 net4290 vdd vss unit_coupling_tile
xi981 net4291 net4088 net4294 net4288 net4287 net4293 net4087 net4292 vdd vss unit_coupling_tile
xi979 net4300 net4093 net4223 net4299 net4296 net4226 net4094 net4295 vdd vss unit_coupling_tile
xi978 net4224 net4096 net4222 net4223 net4226 net4221 net4095 net4225 vdd vss unit_coupling_tile
xi977 net4227 net4020 net4230 net4222 net4221 net4229 net4021 net4228 vdd vss unit_coupling_tile
xi976 net4233 net4023 net4232 net4230 net4229 net4231 net4024 net4234 vdd vss unit_coupling_tile
xi975 net4237 net4029 net4236 net4232 net4231 net4235 net4030 net4238 vdd vss unit_coupling_tile
xi974 net4239 net4033 net4242 net4236 net4235 net4241 net4034 net4240 vdd vss unit_coupling_tile
xi973 net4245 net4035 net4244 net4242 net4241 net4243 net4036 net4246 vdd vss unit_coupling_tile
xi972 net4250 net4041 net4249 net4244 net4243 net4248 net4042 net4247 vdd vss unit_coupling_tile
xi971 net4253 net4046 net4252 net4249 net4248 net4251 net4043 net4254 vdd vss unit_coupling_tile
xi970 net4257 net4049 net4256 net4252 net4251 net4255 net4050 net4258 vdd vss unit_coupling_tile
xi969 net4259 net4053 net4181 net4256 net4255 net4184 net4054 net4260 vdd vss unit_coupling_tile
xi968 net4182 net4055 net4180 net4181 net4184 net4179 net4056 net4183 vdd vss unit_coupling_tile
xi967 net4185 net3978 net4188 net4180 net4179 net4187 net3979 net4186 vdd vss unit_coupling_tile
xi966 net4191 net3981 net4190 net4188 net4187 net4189 net3982 net4192 vdd vss unit_coupling_tile
xi965 net4196 net3987 net4195 net4190 net4189 net4194 net3988 net4193 vdd vss unit_coupling_tile
xi964 net4199 net3992 net4198 net4195 net4194 net4197 net3989 net4200 vdd vss unit_coupling_tile
xi963 net4203 net3995 net4202 net4198 net4197 net4201 net3996 net4204 vdd vss unit_coupling_tile
xi962 net4205 net3999 net4208 net4202 net4201 net4207 net4000 net4206 vdd vss unit_coupling_tile
xi961 net4211 net4001 net4210 net4208 net4207 net4209 net4002 net4212 vdd vss unit_coupling_tile
xi960 net4215 net4007 net4214 net4210 net4209 net4213 net4008 net4216 vdd vss unit_coupling_tile
xi959 net4217 net4011 net4140 net4214 net4213 net4219 net4012 net4218 vdd vss unit_coupling_tile
xi958 net4141 net4013 net4139 net4140 net4219 net4138 net4014 net4220 vdd vss unit_coupling_tile
xi957 net4144 net3937 net4143 net4139 net4138 net4142 net4016 net4145 vdd vss unit_coupling_tile
xi956 net4148 net3940 net4147 net4143 net4142 net4146 net3941 net4149 vdd vss unit_coupling_tile
xi955 net4150 net3944 net4153 net4147 net4146 net4152 net3945 net4151 vdd vss unit_coupling_tile
xi954 net4156 net3946 net4155 net4153 net4152 net4154 net3947 net4157 vdd vss unit_coupling_tile
xi953 net4160 net3952 net4159 net4155 net4154 net4158 net3953 net4161 vdd vss unit_coupling_tile
xi952 net4162 net3956 net4165 net4159 net4158 net4164 net3957 net4163 vdd vss unit_coupling_tile
xi951 net4168 net3958 net4167 net4165 net4164 net4166 net3959 net4169 vdd vss unit_coupling_tile
xi950 net4173 net3964 net4172 net4167 net4166 net4171 net3965 net4170 vdd vss unit_coupling_tile
xi949 net4175 net3969 net4099 net84 net84 net4174 net3966 net4176 vdd vss unit_coupling_tile
xi948 net4177 net3971 net4098 net4099 net4174 net4097 net3972 net4178 vdd vss unit_coupling_tile
xi947 net4102 net3973 net4101 net4098 net4097 net4100 net3974 net4103 vdd vss unit_coupling_tile
xi946 net4106 net3898 net4105 net4101 net4100 net4104 net3899 net4107 vdd vss unit_coupling_tile
xi945 net4108 net3902 net4111 net4105 net4104 net4110 net3903 net4109 vdd vss unit_coupling_tile
xi944 net4114 net3904 net4113 net4111 net4110 net4112 net3905 net4115 vdd vss unit_coupling_tile
xi943 net4119 net3910 net4118 net4113 net4112 net4117 net3911 net4116 vdd vss unit_coupling_tile
xi942 net4122 net3915 net4121 net4118 net4117 net4120 net3912 net4123 vdd vss unit_coupling_tile
xi941 net4126 net3918 net4125 net4121 net4120 net4124 net3919 net4127 vdd vss unit_coupling_tile
xi940 net4128 net3922 net4131 net4125 net4124 net4130 net3923 net4129 vdd vss unit_coupling_tile
xi939 net4134 net3924 net4133 net4131 net4130 net4132 net3925 net4135 vdd vss unit_coupling_tile
xi938 net4136 net3930 net4058 net4133 net4132 net4057 net3931 net4137 vdd vss unit_coupling_tile
xi937 net4061 net3932 net4060 net4058 net4057 net4059 net3933 net4062 vdd vss unit_coupling_tile
xi936 net4066 net3857 net4065 net4060 net4059 net4064 net3858 net4063 vdd vss unit_coupling_tile
xi935 net4069 net3862 net4068 net4065 net4064 net4067 net3859 net4070 vdd vss unit_coupling_tile
xi934 net4073 net3865 net4072 net4068 net4067 net4071 net3866 net4074 vdd vss unit_coupling_tile
xi933 net4075 net3869 net4078 net4072 net4071 net4077 net3870 net4076 vdd vss unit_coupling_tile
xi932 net4081 net3872 net4080 net4078 net4077 net4079 net3871 net4082 vdd vss unit_coupling_tile
xi930 net4084 net3881 net4090 net4083 net4086 net4089 net3882 net4085 vdd vss unit_coupling_tile
xi929 net4093 net3883 net4092 net4090 net4089 net4091 net3884 net4094 vdd vss unit_coupling_tile
xi928 net4096 net3889 net4019 net4092 net4091 net4022 net3890 net4095 vdd vss unit_coupling_tile
xi927 net4020 net3892 net4018 net4019 net4022 net4017 net3891 net4021 vdd vss unit_coupling_tile
xi926 net4023 net3816 net4026 net4018 net4017 net4025 net3817 net4024 vdd vss unit_coupling_tile
xi925 net4029 net3819 net4028 net4026 net4025 net4027 net3820 net4030 vdd vss unit_coupling_tile
xi924 net4033 net3825 net4032 net4028 net4027 net4031 net3826 net4034 vdd vss unit_coupling_tile
xi923 net4035 net3829 net4038 net4032 net4031 net4037 net3830 net4036 vdd vss unit_coupling_tile
xi922 net4041 net3831 net4040 net4038 net4037 net4039 net3832 net4042 vdd vss unit_coupling_tile
xi921 net4046 net3837 net4045 net4040 net4039 net4044 net3838 net4043 vdd vss unit_coupling_tile
xi920 net4049 net3842 net4048 net4045 net4044 net4047 net3839 net4050 vdd vss unit_coupling_tile
xi919 net4053 net3845 net4052 net4048 net4047 net4051 net3846 net4054 vdd vss unit_coupling_tile
xi918 net4055 net3849 net3977 net4052 net4051 net3980 net3850 net4056 vdd vss unit_coupling_tile
xi917 net3978 net3851 net3976 net3977 net3980 net3975 net3852 net3979 vdd vss unit_coupling_tile
xi916 net3981 net3774 net3984 net3976 net3975 net3983 net3775 net3982 vdd vss unit_coupling_tile
xi915 net3987 net3777 net3986 net3984 net3983 net3985 net3778 net3988 vdd vss unit_coupling_tile
xi914 net3992 net3783 net3991 net3986 net3985 net3990 net3784 net3989 vdd vss unit_coupling_tile
xi913 net3995 net3788 net3994 net3991 net3990 net3993 net3785 net3996 vdd vss unit_coupling_tile
xi912 net3999 net3791 net3998 net3994 net3993 net3997 net3792 net4000 vdd vss unit_coupling_tile
xi911 net4001 net3795 net4004 net3998 net3997 net4003 net3796 net4002 vdd vss unit_coupling_tile
xi910 net4007 net3797 net4006 net4004 net4003 net4005 net3798 net4008 vdd vss unit_coupling_tile
xi909 net4011 net3803 net4010 net4006 net4005 net4009 net3804 net4012 vdd vss unit_coupling_tile
xi908 net4013 net3807 net3936 net4010 net4009 net4015 net3808 net4014 vdd vss unit_coupling_tile
xi907 net3937 net3809 net3935 net3936 net4015 net3934 net3810 net4016 vdd vss unit_coupling_tile
xi906 net3940 net3733 net3939 net3935 net3934 net3938 net3812 net3941 vdd vss unit_coupling_tile
xi905 net3944 net3736 net3943 net3939 net3938 net3942 net3737 net3945 vdd vss unit_coupling_tile
xi904 net3946 net3740 net3949 net3943 net3942 net3948 net3741 net3947 vdd vss unit_coupling_tile
xi903 net3952 net3742 net3951 net3949 net3948 net3950 net3743 net3953 vdd vss unit_coupling_tile
xi902 net3956 net3748 net3955 net3951 net3950 net3954 net3749 net3957 vdd vss unit_coupling_tile
xi901 net3958 net3752 net3961 net3955 net3954 net3960 net3753 net3959 vdd vss unit_coupling_tile
xi900 net3964 net3754 net3963 net3961 net3960 net3962 net3755 net3965 vdd vss unit_coupling_tile
xi899 net3969 net3760 net3968 net85 net85 net3967 net3761 net3966 vdd vss unit_coupling_tile
xi898 net3971 net3765 net3895 net3968 net3967 net3970 net3762 net3972 vdd vss unit_coupling_tile
xi897 net3973 net3767 net3894 net3895 net3970 net3893 net3768 net3974 vdd vss unit_coupling_tile
xi896 net3898 net3769 net3897 net3894 net3893 net3896 net3770 net3899 vdd vss unit_coupling_tile
xi895 net3902 net3694 net3901 net3897 net3896 net3900 net3695 net3903 vdd vss unit_coupling_tile
xi894 net3904 net3698 net3907 net3901 net3900 net3906 net3699 net3905 vdd vss unit_coupling_tile
xi893 net3910 net3700 net3909 net3907 net3906 net3908 net3701 net3911 vdd vss unit_coupling_tile
xi892 net3915 net3706 net3914 net3909 net3908 net3913 net3707 net3912 vdd vss unit_coupling_tile
xi891 net3918 net3711 net3917 net3914 net3913 net3916 net3708 net3919 vdd vss unit_coupling_tile
xi890 net3922 net3714 net3921 net3917 net3916 net3920 net3715 net3923 vdd vss unit_coupling_tile
xi889 net3924 net3718 net3927 net3921 net3920 net3926 net3719 net3925 vdd vss unit_coupling_tile
xi888 net3930 net3720 net3929 net3927 net3926 net3928 net3721 net3931 vdd vss unit_coupling_tile
xi887 net3932 net3726 net3854 net3929 net3928 net3853 net3727 net3933 vdd vss unit_coupling_tile
xi886 net3857 net3728 net3856 net3854 net3853 net3855 net3729 net3858 vdd vss unit_coupling_tile
xi885 net3862 net3653 net3861 net3856 net3855 net3860 net3654 net3859 vdd vss unit_coupling_tile
xi884 net3865 net3658 net3864 net3861 net3860 net3863 net3655 net3866 vdd vss unit_coupling_tile
xi883 net3869 net3660 net3868 net3864 net3863 net3867 net3659 net3870 vdd vss unit_coupling_tile
xi881 net3876 net3667 net3874 net3875 net3878 net3873 net3668 net3877 vdd vss unit_coupling_tile
xi880 net3881 net3673 net3880 net3874 net3873 net3879 net3674 net3882 vdd vss unit_coupling_tile
xi879 net3883 net3677 net3886 net3880 net3879 net3885 net3678 net3884 vdd vss unit_coupling_tile
xi878 net3889 net3679 net3888 net3886 net3885 net3887 net3680 net3890 vdd vss unit_coupling_tile
xi877 net3892 net3685 net3815 net3888 net3887 net3818 net3686 net3891 vdd vss unit_coupling_tile
xi876 net3816 net3688 net3814 net3815 net3818 net3813 net3687 net3817 vdd vss unit_coupling_tile
xi875 net3819 net3612 net3822 net3814 net3813 net3821 net3613 net3820 vdd vss unit_coupling_tile
xi874 net3825 net3615 net3824 net3822 net3821 net3823 net3616 net3826 vdd vss unit_coupling_tile
xi873 net3829 net3621 net3828 net3824 net3823 net3827 net3622 net3830 vdd vss unit_coupling_tile
xi872 net3831 net3625 net3834 net3828 net3827 net3833 net3626 net3832 vdd vss unit_coupling_tile
xi871 net3837 net3627 net3836 net3834 net3833 net3835 net3628 net3838 vdd vss unit_coupling_tile
xi870 net3842 net3633 net3841 net3836 net3835 net3840 net3634 net3839 vdd vss unit_coupling_tile
xi869 net3845 net3638 net3844 net3841 net3840 net3843 net3635 net3846 vdd vss unit_coupling_tile
xi868 net3849 net3641 net3848 net3844 net3843 net3847 net3642 net3850 vdd vss unit_coupling_tile
xi867 net3851 net3645 net3773 net3848 net3847 net3776 net3646 net3852 vdd vss unit_coupling_tile
xi866 net3774 net3647 net3772 net3773 net3776 net3771 net3648 net3775 vdd vss unit_coupling_tile
xi865 net3777 net3570 net3780 net3772 net3771 net3779 net3571 net3778 vdd vss unit_coupling_tile
xi864 net3783 net3573 net3782 net3780 net3779 net3781 net3574 net3784 vdd vss unit_coupling_tile
xi863 net3788 net3579 net3787 net3782 net3781 net3786 net3580 net3785 vdd vss unit_coupling_tile
xi862 net3791 net3584 net3790 net3787 net3786 net3789 net3581 net3792 vdd vss unit_coupling_tile
xi861 net3795 net3587 net3794 net3790 net3789 net3793 net3588 net3796 vdd vss unit_coupling_tile
xi860 net3797 net3591 net3800 net3794 net3793 net3799 net3592 net3798 vdd vss unit_coupling_tile
xi859 net3803 net3593 net3802 net3800 net3799 net3801 net3594 net3804 vdd vss unit_coupling_tile
xi858 net3807 net3599 net3806 net3802 net3801 net3805 net3600 net3808 vdd vss unit_coupling_tile
xi857 net3809 net3603 net3732 net3806 net3805 net3811 net3604 net3810 vdd vss unit_coupling_tile
xi856 net3733 net3605 net3731 net3732 net3811 net3730 net3606 net3812 vdd vss unit_coupling_tile
xi855 net3736 net3529 net3735 net3731 net3730 net3734 net3608 net3737 vdd vss unit_coupling_tile
xi854 net3740 net3532 net3739 net3735 net3734 net3738 net3533 net3741 vdd vss unit_coupling_tile
xi853 net3742 net3536 net3745 net3739 net3738 net3744 net3537 net3743 vdd vss unit_coupling_tile
xi852 net3748 net3538 net3747 net3745 net3744 net3746 net3539 net3749 vdd vss unit_coupling_tile
xi851 net3752 net3544 net3751 net3747 net3746 net3750 net3545 net3753 vdd vss unit_coupling_tile
xi850 net3754 net3548 net3757 net3751 net3750 net3756 net3549 net3755 vdd vss unit_coupling_tile
xi849 net3760 net3550 net3759 net86 net86 net3758 net3551 net3761 vdd vss unit_coupling_tile
xi848 net3765 net3556 net3764 net3759 net3758 net3763 net3557 net3762 vdd vss unit_coupling_tile
xi847 net3767 net3561 net3691 net3764 net3763 net3766 net3558 net3768 vdd vss unit_coupling_tile
xi846 net3769 net3563 net3690 net3691 net3766 net3689 net3564 net3770 vdd vss unit_coupling_tile
xi845 net3694 net3565 net3693 net3690 net3689 net3692 net3566 net3695 vdd vss unit_coupling_tile
xi844 net3698 net3490 net3697 net3693 net3692 net3696 net3491 net3699 vdd vss unit_coupling_tile
xi843 net3700 net3494 net3703 net3697 net3696 net3702 net3495 net3701 vdd vss unit_coupling_tile
xi842 net3706 net3496 net3705 net3703 net3702 net3704 net3497 net3707 vdd vss unit_coupling_tile
xi841 net3711 net3502 net3710 net3705 net3704 net3709 net3503 net3708 vdd vss unit_coupling_tile
xi840 net3714 net3507 net3713 net3710 net3709 net3712 net3504 net3715 vdd vss unit_coupling_tile
xi839 net3718 net3510 net3717 net3713 net3712 net3716 net3511 net3719 vdd vss unit_coupling_tile
xi838 net3720 net3514 net3723 net3717 net3716 net3722 net3515 net3721 vdd vss unit_coupling_tile
xi837 net3726 net3516 net3725 net3723 net3722 net3724 net3517 net3727 vdd vss unit_coupling_tile
xi836 net3728 net3522 net3650 net3725 net3724 net3649 net3523 net3729 vdd vss unit_coupling_tile
xi835 net3653 net3524 net3652 net3650 net3649 net3651 net3525 net3654 vdd vss unit_coupling_tile
xi834 net3658 net3450 net3657 net3652 net3651 net3656 net3449 net3655 vdd vss unit_coupling_tile
xi832 net3665 net3457 net3664 net3661 net3662 net3663 net3458 net3666 vdd vss unit_coupling_tile
xi831 net3667 net3461 net3670 net3664 net3663 net3669 net3462 net3668 vdd vss unit_coupling_tile
xi830 net3673 net3463 net3672 net3670 net3669 net3671 net3464 net3674 vdd vss unit_coupling_tile
xi829 net3677 net3469 net3676 net3672 net3671 net3675 net3470 net3678 vdd vss unit_coupling_tile
xi828 net3679 net3473 net3682 net3676 net3675 net3681 net3474 net3680 vdd vss unit_coupling_tile
xi827 net3685 net3475 net3684 net3682 net3681 net3683 net3476 net3686 vdd vss unit_coupling_tile
xi826 net3688 net3481 net3611 net3684 net3683 net3614 net3482 net3687 vdd vss unit_coupling_tile
xi825 net3612 net3484 net3610 net3611 net3614 net3609 net3483 net3613 vdd vss unit_coupling_tile
xi824 net3615 net3408 net3618 net3610 net3609 net3617 net3409 net3616 vdd vss unit_coupling_tile
xi823 net3621 net3411 net3620 net3618 net3617 net3619 net3412 net3622 vdd vss unit_coupling_tile
xi822 net3625 net3417 net3624 net3620 net3619 net3623 net3418 net3626 vdd vss unit_coupling_tile
xi821 net3627 net3421 net3630 net3624 net3623 net3629 net3422 net3628 vdd vss unit_coupling_tile
xi820 net3633 net3423 net3632 net3630 net3629 net3631 net3424 net3634 vdd vss unit_coupling_tile
xi819 net3638 net3429 net3637 net3632 net3631 net3636 net3430 net3635 vdd vss unit_coupling_tile
xi818 net3641 net3434 net3640 net3637 net3636 net3639 net3431 net3642 vdd vss unit_coupling_tile
xi817 net3645 net3437 net3644 net3640 net3639 net3643 net3438 net3646 vdd vss unit_coupling_tile
xi816 net3647 net3441 net3569 net3644 net3643 net3572 net3442 net3648 vdd vss unit_coupling_tile
xi815 net3570 net3443 net3568 net3569 net3572 net3567 net3444 net3571 vdd vss unit_coupling_tile
xi814 net3573 net3366 net3576 net3568 net3567 net3575 net3367 net3574 vdd vss unit_coupling_tile
xi813 net3579 net3369 net3578 net3576 net3575 net3577 net3370 net3580 vdd vss unit_coupling_tile
xi812 net3584 net3375 net3583 net3578 net3577 net3582 net3376 net3581 vdd vss unit_coupling_tile
xi811 net3587 net3380 net3586 net3583 net3582 net3585 net3377 net3588 vdd vss unit_coupling_tile
xi810 net3591 net3383 net3590 net3586 net3585 net3589 net3384 net3592 vdd vss unit_coupling_tile
xi809 net3593 net3387 net3596 net3590 net3589 net3595 net3388 net3594 vdd vss unit_coupling_tile
xi808 net3599 net3389 net3598 net3596 net3595 net3597 net3390 net3600 vdd vss unit_coupling_tile
xi807 net3603 net3395 net3602 net3598 net3597 net3601 net3396 net3604 vdd vss unit_coupling_tile
xi806 net3605 net3399 net3528 net3602 net3601 net3607 net3400 net3606 vdd vss unit_coupling_tile
xi805 net3529 net3401 net3527 net3528 net3607 net3526 net3402 net3608 vdd vss unit_coupling_tile
xi804 net3532 net3325 net3531 net3527 net3526 net3530 net3404 net3533 vdd vss unit_coupling_tile
xi803 net3536 net3328 net3535 net3531 net3530 net3534 net3329 net3537 vdd vss unit_coupling_tile
xi802 net3538 net3332 net3541 net3535 net3534 net3540 net3333 net3539 vdd vss unit_coupling_tile
xi801 net3544 net3334 net3543 net3541 net3540 net3542 net3335 net3545 vdd vss unit_coupling_tile
xi800 net3548 net3340 net3547 net3543 net3542 net3546 net3341 net3549 vdd vss unit_coupling_tile
xi799 net3550 net3344 net3553 net87 net87 net3552 net3345 net3551 vdd vss unit_coupling_tile
xi798 net3556 net3346 net3555 net3553 net3552 net3554 net3347 net3557 vdd vss unit_coupling_tile
xi797 net3561 net3352 net3560 net3555 net3554 net3559 net3353 net3558 vdd vss unit_coupling_tile
xi796 net3563 net3357 net3487 net3560 net3559 net3562 net3354 net3564 vdd vss unit_coupling_tile
xi795 net3565 net3359 net3486 net3487 net3562 net3485 net3360 net3566 vdd vss unit_coupling_tile
xi794 net3490 net3361 net3489 net3486 net3485 net3488 net3362 net3491 vdd vss unit_coupling_tile
xi793 net3494 net3286 net3493 net3489 net3488 net3492 net3287 net3495 vdd vss unit_coupling_tile
xi792 net3496 net3290 net3499 net3493 net3492 net3498 net3291 net3497 vdd vss unit_coupling_tile
xi791 net3502 net3292 net3501 net3499 net3498 net3500 net3293 net3503 vdd vss unit_coupling_tile
xi790 net3507 net3298 net3506 net3501 net3500 net3505 net3299 net3504 vdd vss unit_coupling_tile
xi789 net3510 net3303 net3509 net3506 net3505 net3508 net3300 net3511 vdd vss unit_coupling_tile
xi788 net3514 net3306 net3513 net3509 net3508 net3512 net3307 net3515 vdd vss unit_coupling_tile
xi787 net3516 net3310 net3519 net3513 net3512 net3518 net3311 net3517 vdd vss unit_coupling_tile
xi786 net3522 net3312 net3521 net3519 net3518 net3520 net3313 net3523 vdd vss unit_coupling_tile
xi785 net3524 net3317 net3446 net3521 net3520 net3445 net3316 net3525 vdd vss unit_coupling_tile
xi783 net3454 net3245 net3453 net3451 net3448 net3452 net3246 net3447 vdd vss unit_coupling_tile
xi782 net3457 net3250 net3456 net3453 net3452 net3455 net3247 net3458 vdd vss unit_coupling_tile
xi781 net3461 net3253 net3460 net3456 net3455 net3459 net3254 net3462 vdd vss unit_coupling_tile
xi780 net3463 net3257 net3466 net3460 net3459 net3465 net3258 net3464 vdd vss unit_coupling_tile
xi779 net3469 net3259 net3468 net3466 net3465 net3467 net3260 net3470 vdd vss unit_coupling_tile
xi778 net3473 net3265 net3472 net3468 net3467 net3471 net3266 net3474 vdd vss unit_coupling_tile
xi777 net3475 net3269 net3478 net3472 net3471 net3477 net3270 net3476 vdd vss unit_coupling_tile
xi776 net3481 net3271 net3480 net3478 net3477 net3479 net3272 net3482 vdd vss unit_coupling_tile
xi775 net3484 net3277 net3407 net3480 net3479 net3410 net3278 net3483 vdd vss unit_coupling_tile
xi774 net3408 net3280 net3406 net3407 net3410 net3405 net3279 net3409 vdd vss unit_coupling_tile
xi773 net3411 net3204 net3414 net3406 net3405 net3413 net3205 net3412 vdd vss unit_coupling_tile
xi772 net3417 net3207 net3416 net3414 net3413 net3415 net3208 net3418 vdd vss unit_coupling_tile
xi771 net3421 net3213 net3420 net3416 net3415 net3419 net3214 net3422 vdd vss unit_coupling_tile
xi770 net3423 net3217 net3426 net3420 net3419 net3425 net3218 net3424 vdd vss unit_coupling_tile
xi769 net3429 net3219 net3428 net3426 net3425 net3427 net3220 net3430 vdd vss unit_coupling_tile
xi768 net3434 net3225 net3433 net3428 net3427 net3432 net3226 net3431 vdd vss unit_coupling_tile
xi767 net3437 net3230 net3436 net3433 net3432 net3435 net3227 net3438 vdd vss unit_coupling_tile
xi766 net3441 net3233 net3440 net3436 net3435 net3439 net3234 net3442 vdd vss unit_coupling_tile
xi765 net3443 net3237 net3365 net3440 net3439 net3368 net3238 net3444 vdd vss unit_coupling_tile
xi764 net3366 net3239 net3364 net3365 net3368 net3363 net3240 net3367 vdd vss unit_coupling_tile
xi763 net3369 net3162 net3372 net3364 net3363 net3371 net3163 net3370 vdd vss unit_coupling_tile
xi762 net3375 net3165 net3374 net3372 net3371 net3373 net3166 net3376 vdd vss unit_coupling_tile
xi761 net3380 net3171 net3379 net3374 net3373 net3378 net3172 net3377 vdd vss unit_coupling_tile
xi760 net3383 net3176 net3382 net3379 net3378 net3381 net3173 net3384 vdd vss unit_coupling_tile
xi759 net3387 net3179 net3386 net3382 net3381 net3385 net3180 net3388 vdd vss unit_coupling_tile
xi758 net3389 net3183 net3392 net3386 net3385 net3391 net3184 net3390 vdd vss unit_coupling_tile
xi757 net3395 net3185 net3394 net3392 net3391 net3393 net3186 net3396 vdd vss unit_coupling_tile
xi756 net3399 net3191 net3398 net3394 net3393 net3397 net3192 net3400 vdd vss unit_coupling_tile
xi755 net3401 net3195 net3324 net3398 net3397 net3403 net3196 net3402 vdd vss unit_coupling_tile
xi754 net3325 net3197 net3323 net3324 net3403 net3322 net3198 net3404 vdd vss unit_coupling_tile
xi753 net3328 net3121 net3327 net3323 net3322 net3326 net3200 net3329 vdd vss unit_coupling_tile
xi752 net3332 net3124 net3331 net3327 net3326 net3330 net3125 net3333 vdd vss unit_coupling_tile
xi751 net3334 net3128 net3337 net3331 net3330 net3336 net3129 net3335 vdd vss unit_coupling_tile
xi750 net3340 net3130 net3339 net3337 net3336 net3338 net3131 net3341 vdd vss unit_coupling_tile
xi749 net3344 net3136 net3343 net88 net88 net3342 net3137 net3345 vdd vss unit_coupling_tile
xi748 net3346 net3140 net3349 net3343 net3342 net3348 net3141 net3347 vdd vss unit_coupling_tile
xi747 net3352 net3142 net3351 net3349 net3348 net3350 net3143 net3353 vdd vss unit_coupling_tile
xi746 net3357 net3148 net3356 net3351 net3350 net3355 net3149 net3354 vdd vss unit_coupling_tile
xi745 net3359 net3153 net3283 net3356 net3355 net3358 net3150 net3360 vdd vss unit_coupling_tile
xi744 net3361 net3155 net3282 net3283 net3358 net3281 net3156 net3362 vdd vss unit_coupling_tile
xi743 net3286 net3157 net3285 net3282 net3281 net3284 net3158 net3287 vdd vss unit_coupling_tile
xi742 net3290 net3082 net3289 net3285 net3284 net3288 net3083 net3291 vdd vss unit_coupling_tile
xi741 net3292 net3086 net3295 net3289 net3288 net3294 net3087 net3293 vdd vss unit_coupling_tile
xi740 net3298 net3088 net3297 net3295 net3294 net3296 net3089 net3299 vdd vss unit_coupling_tile
xi739 net3303 net3094 net3302 net3297 net3296 net3301 net3095 net3300 vdd vss unit_coupling_tile
xi738 net3306 net3099 net3305 net3302 net3301 net3304 net3096 net3307 vdd vss unit_coupling_tile
xi737 net3310 net3102 net3309 net3305 net3304 net3308 net3103 net3311 vdd vss unit_coupling_tile
xi736 net3312 net3108 net3315 net3309 net3308 net3314 net3107 net3313 vdd vss unit_coupling_tile
xi734 net3320 net3114 net3242 net3318 net3319 net3241 net3115 net3321 vdd vss unit_coupling_tile
xi733 net3245 net3116 net3244 net3242 net3241 net3243 net3117 net3246 vdd vss unit_coupling_tile
xi732 net3250 net449 net3249 net3244 net3243 net3248 net450 net3247 vdd vss unit_coupling_tile
xi731 net3253 net456 net3252 net3249 net3248 net3251 net451 net3254 vdd vss unit_coupling_tile
xi730 net3257 net461 net3256 net3252 net3251 net3255 net462 net3258 vdd vss unit_coupling_tile
xi729 net3259 net467 net3262 net3256 net3255 net3261 net468 net3260 vdd vss unit_coupling_tile
xi728 net3265 net470 net3264 net3262 net3261 net3263 net471 net3266 vdd vss unit_coupling_tile
xi727 net3269 net479 net3268 net3264 net3263 net3267 net480 net3270 vdd vss unit_coupling_tile
xi726 net3271 net485 net3274 net3268 net3267 net3273 net486 net3272 vdd vss unit_coupling_tile
xi725 net3277 net489 net3276 net3274 net3273 net3275 net490 net3278 vdd vss unit_coupling_tile
xi724 net3280 net497 net3203 net3276 net3275 net3206 net498 net3279 vdd vss unit_coupling_tile
xi723 net3204 net504 net3202 net3203 net3206 net3201 net499 net3205 vdd vss unit_coupling_tile
xi722 net3207 net1183 net3210 net3202 net3201 net3209 net1184 net3208 vdd vss unit_coupling_tile
xi721 net3213 net1186 net3212 net3210 net3209 net3211 net1187 net3214 vdd vss unit_coupling_tile
xi720 net3217 net1195 net3216 net3212 net3211 net3215 net1196 net3218 vdd vss unit_coupling_tile
xi719 net3219 net1201 net3222 net3216 net3215 net3221 net1202 net3220 vdd vss unit_coupling_tile
xi718 net3225 net1205 net3224 net3222 net3221 net3223 net1206 net3226 vdd vss unit_coupling_tile
xi717 net3230 net1213 net3229 net3224 net3223 net3228 net1214 net3227 vdd vss unit_coupling_tile
xi716 net3233 net1220 net3232 net3229 net3228 net3231 net1215 net3234 vdd vss unit_coupling_tile
xi715 net3237 net1225 net3236 net3232 net3231 net3235 net1226 net3238 vdd vss unit_coupling_tile
xi714 net3239 net1231 net3161 net3236 net3235 net3164 net1232 net3240 vdd vss unit_coupling_tile
xi713 net3162 net1234 net3160 net3161 net3164 net3159 net1235 net3163 vdd vss unit_coupling_tile
xi712 net3165 net1020 net3168 net3160 net3159 net3167 net1021 net3166 vdd vss unit_coupling_tile
xi711 net3171 net1025 net3170 net3168 net3167 net3169 net1026 net3172 vdd vss unit_coupling_tile
xi710 net3176 net1033 net3175 net3170 net3169 net3174 net1034 net3173 vdd vss unit_coupling_tile
xi709 net3179 net1040 net3178 net3175 net3174 net3177 net1035 net3180 vdd vss unit_coupling_tile
xi708 net3183 net1045 net3182 net3178 net3177 net3181 net1046 net3184 vdd vss unit_coupling_tile
xi707 net3185 net1051 net3188 net3182 net3181 net3187 net1052 net3186 vdd vss unit_coupling_tile
xi706 net3191 net1054 net3190 net3188 net3187 net3189 net1055 net3192 vdd vss unit_coupling_tile
xi705 net3195 net1063 net3194 net3190 net3189 net3193 net1064 net3196 vdd vss unit_coupling_tile
xi704 net3197 net1069 net3120 net3194 net3193 net3199 net1070 net3198 vdd vss unit_coupling_tile
xi703 net3121 net1073 net3119 net3120 net3199 net3118 net1074 net3200 vdd vss unit_coupling_tile
xi702 net3124 net1082 net3123 net3119 net3118 net3122 net1077 net3125 vdd vss unit_coupling_tile
xi701 net3128 net1087 net3127 net3123 net3122 net3126 net1088 net3129 vdd vss unit_coupling_tile
xi700 net3130 net1093 net3133 net3127 net3126 net3132 net1094 net3131 vdd vss unit_coupling_tile
xi699 net3136 net1096 net3135 net89 net89 net3134 net1097 net3137 vdd vss unit_coupling_tile
xi698 net3140 net1105 net3139 net3135 net3134 net3138 net1106 net3141 vdd vss unit_coupling_tile
xi697 net3142 net1111 net3145 net3139 net3138 net3144 net1112 net3143 vdd vss unit_coupling_tile
xi696 net3148 net1115 net3147 net3145 net3144 net3146 net1116 net3149 vdd vss unit_coupling_tile
xi695 net3153 net1123 net3152 net3147 net3146 net3151 net1124 net3150 vdd vss unit_coupling_tile
xi694 net3155 net1130 net3079 net3152 net3151 net3154 net1125 net3156 vdd vss unit_coupling_tile
xi693 net3157 net1135 net3078 net3079 net3154 net3077 net1136 net3158 vdd vss unit_coupling_tile
xi692 net3082 net1138 net3081 net3078 net3077 net3080 net1139 net3083 vdd vss unit_coupling_tile
xi691 net3086 net1411 net3085 net3081 net3080 net3084 net1412 net3087 vdd vss unit_coupling_tile
xi690 net3088 net1417 net3091 net3085 net3084 net3090 net1418 net3089 vdd vss unit_coupling_tile
xi689 net3094 net1421 net3093 net3091 net3090 net3092 net1422 net3095 vdd vss unit_coupling_tile
xi688 net3099 net1429 net3098 net3093 net3092 net3097 net1430 net3096 vdd vss unit_coupling_tile
xi687 net3102 net1440 net3101 net3098 net3097 net3100 net1431 net3103 vdd vss unit_coupling_tile
xi685 net3104 net1447 net3111 net3109 net3106 net3110 net1448 net3105 vdd vss unit_coupling_tile
xi684 net3114 net1450 net3113 net3111 net3110 net3112 net1451 net3115 vdd vss unit_coupling_tile
xi683 net3116 net1459 net444 net3113 net3112 net443 net1460 net3117 vdd vss unit_coupling_tile
xi682 net449 net447 net446 net444 net443 net445 net448 net450 vdd vss unit_coupling_tile
xi681 net456 net454 net453 net446 net445 net452 net455 net451 vdd vss unit_coupling_tile
xi680 net461 net459 net458 net453 net452 net457 net460 net462 vdd vss unit_coupling_tile
xi679 net467 net465 net464 net458 net457 net463 net466 net468 vdd vss unit_coupling_tile
xi678 net470 net474 net473 net464 net463 net472 net469 net471 vdd vss unit_coupling_tile
xi677 net479 net477 net476 net473 net472 net475 net478 net480 vdd vss unit_coupling_tile
xi676 net485 net483 net482 net476 net475 net481 net484 net486 vdd vss unit_coupling_tile
xi675 net489 net487 net492 net482 net481 net491 net488 net490 vdd vss unit_coupling_tile
xi674 net497 net495 net494 net492 net491 net493 net496 net498 vdd vss unit_coupling_tile
xi673 net504 net502 net501 net494 net493 net500 net503 net499 vdd vss unit_coupling_tile
xi672 net1183 net1181 net1180 net501 net500 net1179 net1182 net1184 vdd vss unit_coupling_tile
xi671 net1186 net1190 net1189 net1180 net1179 net1188 net1185 net1187 vdd vss unit_coupling_tile
xi670 net1195 net1193 net1192 net1189 net1188 net1191 net1194 net1196 vdd vss unit_coupling_tile
xi669 net1201 net1199 net1198 net1192 net1191 net1197 net1200 net1202 vdd vss unit_coupling_tile
xi668 net1205 net1203 net1208 net1198 net1197 net1207 net1204 net1206 vdd vss unit_coupling_tile
xi667 net1213 net1211 net1210 net1208 net1207 net1209 net1212 net1214 vdd vss unit_coupling_tile
xi666 net1220 net1218 net1217 net1210 net1209 net1216 net1219 net1215 vdd vss unit_coupling_tile
xi665 net1225 net1223 net1222 net1217 net1216 net1221 net1224 net1226 vdd vss unit_coupling_tile
xi664 net1231 net1229 net1228 net1222 net1221 net1227 net1230 net1232 vdd vss unit_coupling_tile
xi663 net1234 net1236 net1017 net1228 net1227 net1022 net1233 net1235 vdd vss unit_coupling_tile
xi662 net1020 net1018 net1016 net1017 net1022 net1015 net1019 net1021 vdd vss unit_coupling_tile
xi661 net1025 net1023 net1028 net1016 net1015 net1027 net1024 net1026 vdd vss unit_coupling_tile
xi660 net1033 net1031 net1030 net1028 net1027 net1029 net1032 net1034 vdd vss unit_coupling_tile
xi659 net1040 net1038 net1037 net1030 net1029 net1036 net1039 net1035 vdd vss unit_coupling_tile
xi658 net1045 net1043 net1042 net1037 net1036 net1041 net1044 net1046 vdd vss unit_coupling_tile
xi657 net1051 net1049 net1048 net1042 net1041 net1047 net1050 net1052 vdd vss unit_coupling_tile
xi656 net1054 net1058 net1057 net1048 net1047 net1056 net1053 net1055 vdd vss unit_coupling_tile
xi655 net1063 net1061 net1060 net1057 net1056 net1059 net1062 net1064 vdd vss unit_coupling_tile
xi654 net1069 net1067 net1066 net1060 net1059 net1065 net1068 net1070 vdd vss unit_coupling_tile
xi653 net1073 net1071 net1076 net1066 net1065 net1075 net1072 net1074 vdd vss unit_coupling_tile
xi652 net1082 net1080 net1079 net1076 net1075 net1078 net1081 net1077 vdd vss unit_coupling_tile
xi651 net1087 net1085 net1084 net1079 net1078 net1083 net1086 net1088 vdd vss unit_coupling_tile
xi650 net1093 net1091 net1090 net1084 net1083 net1089 net1092 net1094 vdd vss unit_coupling_tile
xi649 net1096 net1100 net1099 net90 net90 net1098 net1095 net1097 vdd vss unit_coupling_tile
xi648 net1105 net1103 net1102 net1099 net1098 net1101 net1104 net1106 vdd vss unit_coupling_tile
xi647 net1111 net1109 net1108 net1102 net1101 net1107 net1110 net1112 vdd vss unit_coupling_tile
xi646 net1115 net1113 net1118 net1108 net1107 net1117 net1114 net1116 vdd vss unit_coupling_tile
xi645 net1123 net1121 net1120 net1118 net1117 net1119 net1122 net1124 vdd vss unit_coupling_tile
xi644 net1130 net1128 net1127 net1120 net1119 net1126 net1129 net1125 vdd vss unit_coupling_tile
xi643 net1135 net1133 net1132 net1127 net1126 net1131 net1134 net1136 vdd vss unit_coupling_tile
xi642 net1138 net1406 net1405 net1132 net1131 net1404 net1137 net1139 vdd vss unit_coupling_tile
xi641 net1411 net1409 net1408 net1405 net1404 net1407 net1410 net1412 vdd vss unit_coupling_tile
xi640 net1417 net1415 net1414 net1408 net1407 net1413 net1416 net1418 vdd vss unit_coupling_tile
xi639 net1421 net1419 net1424 net1414 net1413 net1423 net1420 net1422 vdd vss unit_coupling_tile
xi638 net1429 net1427 net1426 net1424 net1423 net1425 net1428 net1430 vdd vss unit_coupling_tile
xi636 net1437 net1435 net1433 net1434 net1439 net1432 net1436 net1438 vdd vss unit_coupling_tile
xi635 net1447 net1445 net1444 net1433 net1432 net1443 net1446 net1448 vdd vss unit_coupling_tile
xi634 net1450 net1454 net1453 net1444 net1443 net1452 net1449 net1451 vdd vss unit_coupling_tile
xi633 net1459 net1457 net1456 net1453 net1452 net1455 net1458 net1460 vdd vss unit_coupling_tile
xi632 net447 net1461 net1260 net1456 net1455 net1259 net1462 net448 vdd vss unit_coupling_tile
xi631 net454 net1263 net1262 net1260 net1259 net1261 net1264 net455 vdd vss unit_coupling_tile
xi630 net459 net1267 net1266 net1262 net1261 net1265 net1268 net460 vdd vss unit_coupling_tile
xi629 net465 net1271 net1270 net1266 net1265 net1269 net1272 net466 vdd vss unit_coupling_tile
xi628 net474 net1275 net1274 net1270 net1269 net1273 net1276 net469 vdd vss unit_coupling_tile
xi627 net477 net1280 net1279 net1274 net1273 net1278 net1277 net478 vdd vss unit_coupling_tile
xi626 net483 net1283 net1282 net1279 net1278 net1281 net1284 net484 vdd vss unit_coupling_tile
xi625 net487 net1287 net1286 net1282 net1281 net1285 net1288 net488 vdd vss unit_coupling_tile
xi624 net495 net1289 net1292 net1286 net1285 net1291 net1290 net496 vdd vss unit_coupling_tile
xi623 net502 net1295 net1294 net1292 net1291 net1293 net1296 net503 vdd vss unit_coupling_tile
xi622 net1181 net1299 net1298 net1294 net1293 net1297 net1300 net1182 vdd vss unit_coupling_tile
xi621 net1190 net1368 net1367 net1298 net1297 net1366 net1369 net1185 vdd vss unit_coupling_tile
xi620 net1193 net1373 net1372 net1367 net1366 net1371 net1370 net1194 vdd vss unit_coupling_tile
xi619 net1199 net1376 net1375 net1372 net1371 net1374 net1377 net1200 vdd vss unit_coupling_tile
xi618 net1203 net1380 net1379 net1375 net1374 net1378 net1381 net1204 vdd vss unit_coupling_tile
xi617 net1211 net1382 net1385 net1379 net1378 net1384 net1383 net1212 vdd vss unit_coupling_tile
xi616 net1218 net1388 net1387 net1385 net1384 net1386 net1389 net1219 vdd vss unit_coupling_tile
xi615 net1223 net1392 net1391 net1387 net1386 net1390 net1393 net1224 vdd vss unit_coupling_tile
xi614 net1229 net1396 net1395 net1391 net1390 net1394 net1397 net1230 vdd vss unit_coupling_tile
xi613 net1236 net1400 net1399 net1395 net1394 net1398 net1401 net1233 vdd vss unit_coupling_tile
xi612 net1018 net1403 net1303 net1399 net1398 net1306 net1402 net1019 vdd vss unit_coupling_tile
xi611 net1023 net1304 net1302 net1303 net1306 net1301 net1305 net1024 vdd vss unit_coupling_tile
xi610 net1031 net1307 net1310 net1302 net1301 net1309 net1308 net1032 vdd vss unit_coupling_tile
xi609 net1038 net1313 net1312 net1310 net1309 net1311 net1314 net1039 vdd vss unit_coupling_tile
xi608 net1043 net1317 net1316 net1312 net1311 net1315 net1318 net1044 vdd vss unit_coupling_tile
xi607 net1049 net1321 net1320 net1316 net1315 net1319 net1322 net1050 vdd vss unit_coupling_tile
xi606 net1058 net1325 net1324 net1320 net1319 net1323 net1326 net1053 vdd vss unit_coupling_tile
xi605 net1061 net1330 net1329 net1324 net1323 net1328 net1327 net1062 vdd vss unit_coupling_tile
xi604 net1067 net1333 net1332 net1329 net1328 net1331 net1334 net1068 vdd vss unit_coupling_tile
xi603 net1071 net1337 net1336 net1332 net1331 net1335 net1338 net1072 vdd vss unit_coupling_tile
xi602 net1080 net1339 net1342 net1336 net1335 net1341 net1340 net1081 vdd vss unit_coupling_tile
xi601 net1085 net1543 net1835 net1342 net1341 net1834 net1544 net1086 vdd vss unit_coupling_tile
xi600 net1091 net1654 net1837 net1835 net1834 net1836 net1547 net1092 vdd vss unit_coupling_tile
xi599 net1100 net1659 net1839 net91 net91 net1838 net1660 net1095 vdd vss unit_coupling_tile
xi598 net1103 net1665 net1841 net1839 net1838 net1840 net1666 net1104 vdd vss unit_coupling_tile
xi597 net1109 net1668 net1843 net1841 net1840 net1842 net1669 net1110 vdd vss unit_coupling_tile
xi596 net1113 net1677 net1845 net1843 net1842 net1844 net1678 net1114 vdd vss unit_coupling_tile
xi595 net1121 net1683 net1847 net1845 net1844 net1846 net1684 net1122 vdd vss unit_coupling_tile
xi594 net1128 net1687 net1849 net1847 net1846 net1848 net1688 net1129 vdd vss unit_coupling_tile
xi593 net1133 net1695 net1851 net1849 net1848 net1850 net1696 net1134 vdd vss unit_coupling_tile
xi592 net1406 net1702 net1853 net1851 net1850 net1852 net1697 net1137 vdd vss unit_coupling_tile
xi591 net1409 net1707 net1855 net1853 net1852 net1854 net1708 net1410 vdd vss unit_coupling_tile
xi590 net1415 net1710 net1857 net1855 net1854 net1856 net1711 net1416 vdd vss unit_coupling_tile
xi589 net1419 net1716 net1859 net1857 net1856 net1858 net1715 net1420 vdd vss unit_coupling_tile
xi587 net1442 net1729 net1861 net1862 net1863 net1860 net1730 net1441 vdd vss unit_coupling_tile
xi586 net1435 net1737 net1865 net1861 net1860 net1864 net1738 net1436 vdd vss unit_coupling_tile
xi585 net1445 net1744 net1867 net1865 net1864 net1866 net1739 net1446 vdd vss unit_coupling_tile
xi584 net1454 net1749 net1869 net1867 net1866 net1868 net1750 net1449 vdd vss unit_coupling_tile
xi583 net1457 net1755 net1871 net1869 net1868 net1870 net1756 net1458 vdd vss unit_coupling_tile
xi582 net1461 net1758 net1873 net1871 net1870 net1872 net1759 net1462 vdd vss unit_coupling_tile
xi581 net1263 net1767 net1875 net1873 net1872 net1874 net1768 net1264 vdd vss unit_coupling_tile
xi580 net1267 net1771 net1877 net1875 net1874 net1876 net1772 net1268 vdd vss unit_coupling_tile
xi579 net1271 net1598 net1879 net1877 net1876 net1878 net1599 net1272 vdd vss unit_coupling_tile
xi578 net1275 net1605 net1881 net1879 net1878 net1880 net1600 net1276 vdd vss unit_coupling_tile
xi577 net1280 net1610 net1883 net1881 net1880 net1882 net1611 net1277 vdd vss unit_coupling_tile
xi576 net1283 net1616 net1885 net1883 net1882 net1884 net1617 net1284 vdd vss unit_coupling_tile
xi575 net1287 net1619 net1887 net1885 net1884 net1886 net1620 net1288 vdd vss unit_coupling_tile
xi574 net1289 net1628 net1889 net1887 net1886 net1888 net1629 net1290 vdd vss unit_coupling_tile
xi573 net1295 net1634 net1891 net1889 net1888 net1890 net1635 net1296 vdd vss unit_coupling_tile
xi572 net1299 net1638 net1893 net1891 net1890 net1892 net1639 net1300 vdd vss unit_coupling_tile
xi571 net1368 net1646 net1465 net1893 net1892 net1468 net1647 net1369 vdd vss unit_coupling_tile
xi570 net1373 net1466 net1464 net1465 net1468 net1463 net1467 net1370 vdd vss unit_coupling_tile
xi569 net1376 net1472 net1471 net1464 net1463 net1470 net1469 net1377 vdd vss unit_coupling_tile
xi568 net1380 net1475 net1474 net1471 net1470 net1473 net1476 net1381 vdd vss unit_coupling_tile
xi567 net1382 net1479 net1478 net1474 net1473 net1477 net1480 net1383 vdd vss unit_coupling_tile
xi566 net1388 net1481 net1484 net1478 net1477 net1483 net1482 net1389 vdd vss unit_coupling_tile
xi565 net1392 net1487 net1486 net1484 net1483 net1485 net1488 net1393 vdd vss unit_coupling_tile
xi564 net1396 net1491 net1490 net1486 net1485 net1489 net1492 net1397 vdd vss unit_coupling_tile
xi563 net1400 net1495 net1494 net1490 net1489 net1493 net1496 net1401 vdd vss unit_coupling_tile
xi562 net1403 net1499 net1498 net1494 net1493 net1497 net1500 net1402 vdd vss unit_coupling_tile
xi561 net1304 net1504 net1503 net1498 net1497 net1502 net1501 net1305 vdd vss unit_coupling_tile
xi560 net1307 net1507 net1506 net1503 net1502 net1505 net1508 net1308 vdd vss unit_coupling_tile
xi559 net1313 net1509 net1512 net1506 net1505 net1511 net1510 net1314 vdd vss unit_coupling_tile
xi558 net1317 net1515 net1514 net1512 net1511 net1513 net1516 net1318 vdd vss unit_coupling_tile
xi557 net1321 net1519 net1518 net1514 net1513 net1517 net1520 net1322 vdd vss unit_coupling_tile
xi556 net1325 net1523 net1522 net1518 net1517 net1521 net1524 net1326 vdd vss unit_coupling_tile
xi555 net1330 net1527 net1526 net1522 net1521 net1525 net1528 net1327 vdd vss unit_coupling_tile
xi554 net1333 net1532 net1531 net1526 net1525 net1530 net1529 net1334 vdd vss unit_coupling_tile
xi553 net1337 net1535 net1534 net1531 net1530 net1533 net1536 net1338 vdd vss unit_coupling_tile
xi552 net1339 net1539 net1538 net1534 net1533 net1537 net1540 net1340 vdd vss unit_coupling_tile
xi551 net1543 net1541 net1546 net1538 net1537 net1545 net1542 net1544 vdd vss unit_coupling_tile
xi550 net1654 net1652 net1651 net1546 net1545 net1650 net1653 net1547 vdd vss unit_coupling_tile
xi549 net1659 net1657 net1656 net92 net92 net1655 net1658 net1660 vdd vss unit_coupling_tile
xi548 net1665 net1663 net1662 net1656 net1655 net1661 net1664 net1666 vdd vss unit_coupling_tile
xi547 net1668 net1672 net1671 net1662 net1661 net1670 net1667 net1669 vdd vss unit_coupling_tile
xi546 net1677 net1675 net1674 net1671 net1670 net1673 net1676 net1678 vdd vss unit_coupling_tile
xi545 net1683 net1681 net1680 net1674 net1673 net1679 net1682 net1684 vdd vss unit_coupling_tile
xi544 net1687 net1685 net1690 net1680 net1679 net1689 net1686 net1688 vdd vss unit_coupling_tile
xi543 net1695 net1693 net1692 net1690 net1689 net1691 net1694 net1696 vdd vss unit_coupling_tile
xi542 net1702 net1700 net1699 net1692 net1691 net1698 net1701 net1697 vdd vss unit_coupling_tile
xi541 net1707 net1705 net1704 net1699 net1698 net1703 net1706 net1708 vdd vss unit_coupling_tile
xi540 net1710 net1714 net1713 net1704 net1703 net1712 net1709 net1711 vdd vss unit_coupling_tile
xi538 net1725 net1723 net1722 net1719 net1720 net1721 net1724 net1726 vdd vss unit_coupling_tile
xi537 net1729 net1727 net1732 net1722 net1721 net1731 net1728 net1730 vdd vss unit_coupling_tile
xi536 net1737 net1735 net1734 net1732 net1731 net1733 net1736 net1738 vdd vss unit_coupling_tile
xi535 net1744 net1742 net1741 net1734 net1733 net1740 net1743 net1739 vdd vss unit_coupling_tile
xi534 net1749 net1747 net1746 net1741 net1740 net1745 net1748 net1750 vdd vss unit_coupling_tile
xi533 net1755 net1753 net1752 net1746 net1745 net1751 net1754 net1756 vdd vss unit_coupling_tile
xi532 net1758 net1762 net1761 net1752 net1751 net1760 net1757 net1759 vdd vss unit_coupling_tile
xi531 net1767 net1765 net1764 net1761 net1760 net1763 net1766 net1768 vdd vss unit_coupling_tile
xi530 net1771 net1769 net1593 net1764 net1763 net1592 net1770 net1772 vdd vss unit_coupling_tile
xi529 net1598 net1596 net1595 net1593 net1592 net1594 net1597 net1599 vdd vss unit_coupling_tile
xi528 net1605 net1603 net1602 net1595 net1594 net1601 net1604 net1600 vdd vss unit_coupling_tile
xi527 net1610 net1608 net1607 net1602 net1601 net1606 net1609 net1611 vdd vss unit_coupling_tile
xi526 net1616 net1614 net1613 net1607 net1606 net1612 net1615 net1617 vdd vss unit_coupling_tile
xi525 net1619 net1623 net1622 net1613 net1612 net1621 net1618 net1620 vdd vss unit_coupling_tile
xi524 net1628 net1626 net1625 net1622 net1621 net1624 net1627 net1629 vdd vss unit_coupling_tile
xi523 net1634 net1632 net1631 net1625 net1624 net1630 net1633 net1635 vdd vss unit_coupling_tile
xi522 net1638 net1636 net1641 net1631 net1630 net1640 net1637 net1639 vdd vss unit_coupling_tile
xi521 net1646 net1644 net1643 net1641 net1640 net1642 net1645 net1647 vdd vss unit_coupling_tile
xi520 net1466 net1648 net1550 net1643 net1642 net1553 net1649 net1467 vdd vss unit_coupling_tile
xi519 net1472 net1551 net1549 net1550 net1553 net1548 net1552 net1469 vdd vss unit_coupling_tile
xi518 net1475 net1557 net1556 net1549 net1548 net1555 net1554 net1476 vdd vss unit_coupling_tile
xi517 net1479 net1560 net1559 net1556 net1555 net1558 net1561 net1480 vdd vss unit_coupling_tile
xi516 net1481 net1564 net1563 net1559 net1558 net1562 net1565 net1482 vdd vss unit_coupling_tile
xi515 net1487 net1566 net1569 net1563 net1562 net1568 net1567 net1488 vdd vss unit_coupling_tile
xi514 net1491 net1572 net1571 net1569 net1568 net1570 net1573 net1492 vdd vss unit_coupling_tile
xi513 net1495 net1576 net1575 net1571 net1570 net1574 net1577 net1496 vdd vss unit_coupling_tile
xi512 net1499 net1580 net1579 net1575 net1574 net1578 net1581 net1500 vdd vss unit_coupling_tile
xi511 net1504 net1584 net1583 net1579 net1578 net1582 net1585 net1501 vdd vss unit_coupling_tile
xi510 net1507 net1589 net1588 net1583 net1582 net1587 net1586 net1508 vdd vss unit_coupling_tile
xi509 net1509 net1915 net1914 net1588 net1587 net1913 net1916 net1510 vdd vss unit_coupling_tile
xi508 net1515 net1917 net1920 net1914 net1913 net1919 net1918 net1516 vdd vss unit_coupling_tile
xi507 net1519 net1923 net1922 net1920 net1919 net1921 net1924 net1520 vdd vss unit_coupling_tile
xi506 net1523 net1927 net1926 net1922 net1921 net1925 net1928 net1524 vdd vss unit_coupling_tile
xi505 net1527 net1931 net1930 net1926 net1925 net1929 net1932 net1528 vdd vss unit_coupling_tile
xi504 net1532 net1935 net1934 net1930 net1929 net1933 net1936 net1529 vdd vss unit_coupling_tile
xi503 net1535 net1940 net1939 net1934 net1933 net1938 net1937 net1536 vdd vss unit_coupling_tile
xi502 net1539 net1943 net1942 net1939 net1938 net1941 net1944 net1540 vdd vss unit_coupling_tile
xi501 net1541 net1947 net1946 net1942 net1941 net1945 net1948 net1542 vdd vss unit_coupling_tile
xi500 net1652 net1949 net1952 net1946 net1945 net1951 net1950 net1653 vdd vss unit_coupling_tile
xi499 net1657 net1955 net1954 net93 net93 net1953 net1956 net1658 vdd vss unit_coupling_tile
xi498 net1663 net1959 net1958 net1954 net1953 net1957 net1960 net1664 vdd vss unit_coupling_tile
xi497 net1672 net1963 net1962 net1958 net1957 net1961 net1964 net1667 vdd vss unit_coupling_tile
xi496 net1675 net1968 net1967 net1962 net1961 net1966 net1965 net1676 vdd vss unit_coupling_tile
xi495 net1681 net1971 net1970 net1967 net1966 net1969 net1972 net1682 vdd vss unit_coupling_tile
xi494 net1685 net1975 net1974 net1970 net1969 net1973 net1976 net1686 vdd vss unit_coupling_tile
xi493 net1693 net1977 net1980 net1974 net1973 net1979 net1978 net1694 vdd vss unit_coupling_tile
xi492 net1700 net1983 net1982 net1980 net1979 net1981 net1984 net1701 vdd vss unit_coupling_tile
xi491 net1705 net1987 net1986 net1982 net1981 net1985 net1988 net1706 vdd vss unit_coupling_tile
xi489 net1718 net1996 net1995 net1991 net1992 net1994 net1993 net1717 vdd vss unit_coupling_tile
xi488 net1723 net1999 net1998 net1995 net1994 net1997 net2000 net1724 vdd vss unit_coupling_tile
xi487 net1727 net2003 net2002 net1998 net1997 net2001 net2004 net1728 vdd vss unit_coupling_tile
xi486 net1735 net2005 net2008 net2002 net2001 net2007 net2006 net1736 vdd vss unit_coupling_tile
xi485 net1742 net2011 net2010 net2008 net2007 net2009 net2012 net1743 vdd vss unit_coupling_tile
xi484 net1747 net2015 net2014 net2010 net2009 net2013 net2016 net1748 vdd vss unit_coupling_tile
xi483 net1753 net2019 net2018 net2014 net2013 net2017 net2020 net1754 vdd vss unit_coupling_tile
xi482 net1762 net2023 net2022 net2018 net2017 net2021 net2024 net1757 vdd vss unit_coupling_tile
xi481 net1765 net2028 net2027 net2022 net2021 net2026 net2025 net1766 vdd vss unit_coupling_tile
xi480 net1769 net2031 net2030 net2027 net2026 net2029 net2032 net1770 vdd vss unit_coupling_tile
xi479 net1596 net2033 net2036 net2030 net2029 net2035 net2034 net1597 vdd vss unit_coupling_tile
xi478 net1603 net2039 net2038 net2036 net2035 net2037 net2040 net1604 vdd vss unit_coupling_tile
xi477 net1608 net2043 net2042 net2038 net2037 net2041 net2044 net1609 vdd vss unit_coupling_tile
xi476 net1614 net2047 net2046 net2042 net2041 net2045 net2048 net1615 vdd vss unit_coupling_tile
xi475 net1623 net2051 net2050 net2046 net2045 net2049 net2052 net1618 vdd vss unit_coupling_tile
xi474 net1626 net2056 net2055 net2050 net2049 net2054 net2053 net1627 vdd vss unit_coupling_tile
xi473 net1632 net2059 net2058 net2055 net2054 net2057 net2060 net1633 vdd vss unit_coupling_tile
xi472 net1636 net2063 net2062 net2058 net2057 net2061 net2064 net1637 vdd vss unit_coupling_tile
xi471 net1644 net2065 net2068 net2062 net2061 net2067 net2066 net1645 vdd vss unit_coupling_tile
xi470 net1648 net2071 net2070 net2068 net2067 net2069 net2072 net1649 vdd vss unit_coupling_tile
xi469 net1551 net2075 net2074 net2070 net2069 net2073 net2076 net1552 vdd vss unit_coupling_tile
xi468 net1557 net2079 net2078 net2074 net2073 net2077 net2080 net1554 vdd vss unit_coupling_tile
xi467 net1560 net2084 net2083 net2078 net2077 net2082 net2081 net1561 vdd vss unit_coupling_tile
xi466 net1564 net2087 net2086 net2083 net2082 net2085 net2088 net1565 vdd vss unit_coupling_tile
xi465 net1566 net2091 net2090 net2086 net2085 net2089 net2092 net1567 vdd vss unit_coupling_tile
xi464 net1572 net2093 net2096 net2090 net2089 net2095 net2094 net1573 vdd vss unit_coupling_tile
xi463 net1576 net2099 net2098 net2096 net2095 net2097 net2100 net1577 vdd vss unit_coupling_tile
xi462 net1580 net2103 net2102 net2098 net2097 net2101 net2104 net1581 vdd vss unit_coupling_tile
xi461 net1584 net2107 net2106 net2102 net2101 net2105 net2108 net1585 vdd vss unit_coupling_tile
xi460 net1589 net2111 net2110 net2106 net2105 net2109 net2112 net1586 vdd vss unit_coupling_tile
xi459 net1915 net2116 net2115 net2110 net2109 net2114 net2113 net1916 vdd vss unit_coupling_tile
xi458 net1917 net2119 net2118 net2115 net2114 net2117 net2120 net1918 vdd vss unit_coupling_tile
xi457 net1923 net2121 net2124 net2118 net2117 net2123 net2122 net1924 vdd vss unit_coupling_tile
xi456 net1927 net2127 net2126 net2124 net2123 net2125 net2128 net1928 vdd vss unit_coupling_tile
xi455 net1931 net2131 net2130 net2126 net2125 net2129 net2132 net1932 vdd vss unit_coupling_tile
xi454 net1935 net2135 net2134 net2130 net2129 net2133 net2136 net1936 vdd vss unit_coupling_tile
xi453 net1940 net2139 net2138 net2134 net2133 net2137 net2140 net1937 vdd vss unit_coupling_tile
xi452 net1943 net2144 net2143 net2138 net2137 net2142 net2141 net1944 vdd vss unit_coupling_tile
xi451 net1947 net2147 net2146 net2143 net2142 net2145 net2148 net1948 vdd vss unit_coupling_tile
xi450 net1949 net2151 net2150 net2146 net2145 net2149 net2152 net1950 vdd vss unit_coupling_tile
xi449 net1955 net2153 net2156 net94 net94 net2155 net2154 net1956 vdd vss unit_coupling_tile
xi448 net1959 net2159 net2158 net2156 net2155 net2157 net2160 net1960 vdd vss unit_coupling_tile
xi447 net1963 net2163 net2162 net2158 net2157 net2161 net2164 net1964 vdd vss unit_coupling_tile
xi446 net1968 net2167 net2166 net2162 net2161 net2165 net2168 net1965 vdd vss unit_coupling_tile
xi445 net1971 net2172 net2171 net2166 net2165 net2170 net2169 net1972 vdd vss unit_coupling_tile
xi444 net1975 net2175 net2174 net2171 net2170 net2173 net2176 net1976 vdd vss unit_coupling_tile
xi443 net1977 net2179 net2178 net2174 net2173 net2177 net2180 net1978 vdd vss unit_coupling_tile
xi442 net1983 net2181 net2184 net2178 net2177 net2183 net2182 net1984 vdd vss unit_coupling_tile
xi440 net1990 net2191 net2190 net2188 net2185 net2189 net2192 net1989 vdd vss unit_coupling_tile
xi439 net1996 net2195 net2194 net2190 net2189 net2193 net2196 net1993 vdd vss unit_coupling_tile
xi438 net1999 net2200 net2199 net2194 net2193 net2198 net2197 net2000 vdd vss unit_coupling_tile
xi437 net2003 net2203 net2202 net2199 net2198 net2201 net2204 net2004 vdd vss unit_coupling_tile
xi436 net2005 net2207 net2206 net2202 net2201 net2205 net2208 net2006 vdd vss unit_coupling_tile
xi435 net2011 net2209 net2212 net2206 net2205 net2211 net2210 net2012 vdd vss unit_coupling_tile
xi434 net2015 net2215 net2214 net2212 net2211 net2213 net2216 net2016 vdd vss unit_coupling_tile
xi433 net2019 net2219 net2218 net2214 net2213 net2217 net2220 net2020 vdd vss unit_coupling_tile
xi432 net2023 net2223 net2222 net2218 net2217 net2221 net2224 net2024 vdd vss unit_coupling_tile
xi431 net2028 net2227 net2226 net2222 net2221 net2225 net2228 net2025 vdd vss unit_coupling_tile
xi430 net2031 net2232 net2231 net2226 net2225 net2230 net2229 net2032 vdd vss unit_coupling_tile
xi429 net2033 net2235 net2234 net2231 net2230 net2233 net2236 net2034 vdd vss unit_coupling_tile
xi428 net2039 net2237 net2240 net2234 net2233 net2239 net2238 net2040 vdd vss unit_coupling_tile
xi427 net2043 net2243 net2242 net2240 net2239 net2241 net2244 net2044 vdd vss unit_coupling_tile
xi426 net2047 net2247 net2246 net2242 net2241 net2245 net2248 net2048 vdd vss unit_coupling_tile
xi425 net2051 net2251 net2250 net2246 net2245 net2249 net2252 net2052 vdd vss unit_coupling_tile
xi424 net2056 net2255 net2254 net2250 net2249 net2253 net2256 net2053 vdd vss unit_coupling_tile
xi423 net2059 net2260 net2259 net2254 net2253 net2258 net2257 net2060 vdd vss unit_coupling_tile
xi422 net2063 net2263 net2262 net2259 net2258 net2261 net2264 net2064 vdd vss unit_coupling_tile
xi421 net2065 net2267 net2266 net2262 net2261 net2265 net2268 net2066 vdd vss unit_coupling_tile
xi420 net2071 net2269 net2272 net2266 net2265 net2271 net2270 net2072 vdd vss unit_coupling_tile
xi419 net2075 net2275 net2274 net2272 net2271 net2273 net2276 net2076 vdd vss unit_coupling_tile
xi418 net2079 net2279 net2278 net2274 net2273 net2277 net2280 net2080 vdd vss unit_coupling_tile
xi417 net2084 net2283 net2282 net2278 net2277 net2281 net2284 net2081 vdd vss unit_coupling_tile
xi416 net2087 net2288 net2287 net2282 net2281 net2286 net2285 net2088 vdd vss unit_coupling_tile
xi415 net2091 net2291 net2290 net2287 net2286 net2289 net2292 net2092 vdd vss unit_coupling_tile
xi414 net2093 net2295 net2294 net2290 net2289 net2293 net2296 net2094 vdd vss unit_coupling_tile
xi413 net2099 net2297 net2300 net2294 net2293 net2299 net2298 net2100 vdd vss unit_coupling_tile
xi412 net2103 net2303 net2302 net2300 net2299 net2301 net2304 net2104 vdd vss unit_coupling_tile
xi411 net2107 net2307 net2306 net2302 net2301 net2305 net2308 net2108 vdd vss unit_coupling_tile
xi410 net2111 net2311 net2310 net2306 net2305 net2309 net2312 net2112 vdd vss unit_coupling_tile
xi409 net2116 net2315 net2314 net2310 net2309 net2313 net2316 net2113 vdd vss unit_coupling_tile
xi408 net2119 net2320 net2319 net2314 net2313 net2318 net2317 net2120 vdd vss unit_coupling_tile
xi407 net2121 net2323 net2322 net2319 net2318 net2321 net2324 net2122 vdd vss unit_coupling_tile
xi406 net2127 net2325 net2328 net2322 net2321 net2327 net2326 net2128 vdd vss unit_coupling_tile
xi405 net2131 net2331 net2330 net2328 net2327 net2329 net2332 net2132 vdd vss unit_coupling_tile
xi404 net2135 net2335 net2334 net2330 net2329 net2333 net2336 net2136 vdd vss unit_coupling_tile
xi403 net2139 net2339 net2338 net2334 net2333 net2337 net2340 net2140 vdd vss unit_coupling_tile
xi402 net2144 net2343 net2342 net2338 net2337 net2341 net2344 net2141 vdd vss unit_coupling_tile
xi401 net2147 net2348 net2347 net2342 net2341 net2346 net2345 net2148 vdd vss unit_coupling_tile
xi400 net2151 net2351 net2350 net2347 net2346 net2349 net2352 net2152 vdd vss unit_coupling_tile
xi399 net2153 net2355 net2354 net95 net95 net2353 net2356 net2154 vdd vss unit_coupling_tile
xi398 net2159 net2357 net2360 net2354 net2353 net2359 net2358 net2160 vdd vss unit_coupling_tile
xi397 net2163 net2363 net2362 net2360 net2359 net2361 net2364 net2164 vdd vss unit_coupling_tile
xi396 net2167 net2367 net2366 net2362 net2361 net2365 net2368 net2168 vdd vss unit_coupling_tile
xi395 net2172 net2371 net2370 net2366 net2365 net2369 net2372 net2169 vdd vss unit_coupling_tile
xi394 net2175 net2376 net2375 net2370 net2369 net2374 net2373 net2176 vdd vss unit_coupling_tile
xi393 net2179 net2379 net2378 net2375 net2374 net2377 net2380 net2180 vdd vss unit_coupling_tile
xi391 net2187 net2382 net2388 net2381 net2384 net2387 net2383 net2186 vdd vss unit_coupling_tile
xi390 net2191 net2391 net2390 net2388 net2387 net2389 net2392 net2192 vdd vss unit_coupling_tile
xi389 net2195 net2395 net2394 net2390 net2389 net2393 net2396 net2196 vdd vss unit_coupling_tile
xi388 net2200 net2399 net2398 net2394 net2393 net2397 net2400 net2197 vdd vss unit_coupling_tile
xi387 net2203 net2404 net2403 net2398 net2397 net2402 net2401 net2204 vdd vss unit_coupling_tile
xi386 net2207 net2407 net2406 net2403 net2402 net2405 net2408 net2208 vdd vss unit_coupling_tile
xi385 net2209 net2411 net2410 net2406 net2405 net2409 net2412 net2210 vdd vss unit_coupling_tile
xi384 net2215 net2413 net2416 net2410 net2409 net2415 net2414 net2216 vdd vss unit_coupling_tile
xi383 net2219 net2419 net2418 net2416 net2415 net2417 net2420 net2220 vdd vss unit_coupling_tile
xi382 net2223 net2423 net2422 net2418 net2417 net2421 net2424 net2224 vdd vss unit_coupling_tile
xi381 net2227 net2427 net2426 net2422 net2421 net2425 net2428 net2228 vdd vss unit_coupling_tile
xi380 net2232 net2431 net2430 net2426 net2425 net2429 net2432 net2229 vdd vss unit_coupling_tile
xi379 net2235 net2436 net2435 net2430 net2429 net2434 net2433 net2236 vdd vss unit_coupling_tile
xi378 net2237 net2439 net2438 net2435 net2434 net2437 net2440 net2238 vdd vss unit_coupling_tile
xi377 net2243 net2441 net2444 net2438 net2437 net2443 net2442 net2244 vdd vss unit_coupling_tile
xi376 net2247 net2447 net2446 net2444 net2443 net2445 net2448 net2248 vdd vss unit_coupling_tile
xi375 net2251 net2451 net2450 net2446 net2445 net2449 net2452 net2252 vdd vss unit_coupling_tile
xi374 net2255 net2455 net2454 net2450 net2449 net2453 net2456 net2256 vdd vss unit_coupling_tile
xi373 net2260 net2459 net2458 net2454 net2453 net2457 net2460 net2257 vdd vss unit_coupling_tile
xi372 net2263 net2464 net2463 net2458 net2457 net2462 net2461 net2264 vdd vss unit_coupling_tile
xi371 net2267 net2467 net2466 net2463 net2462 net2465 net2468 net2268 vdd vss unit_coupling_tile
xi370 net2269 net2471 net2470 net2466 net2465 net2469 net2472 net2270 vdd vss unit_coupling_tile
xi369 net2275 net2473 net2476 net2470 net2469 net2475 net2474 net2276 vdd vss unit_coupling_tile
xi368 net2279 net2479 net2478 net2476 net2475 net2477 net2480 net2280 vdd vss unit_coupling_tile
xi367 net2283 net2483 net2482 net2478 net2477 net2481 net2484 net2284 vdd vss unit_coupling_tile
xi366 net2288 net2487 net2486 net2482 net2481 net2485 net2488 net2285 vdd vss unit_coupling_tile
xi365 net2291 net2492 net2491 net2486 net2485 net2490 net2489 net2292 vdd vss unit_coupling_tile
xi364 net2295 net2495 net2494 net2491 net2490 net2493 net2496 net2296 vdd vss unit_coupling_tile
xi363 net2297 net2499 net2498 net2494 net2493 net2497 net2500 net2298 vdd vss unit_coupling_tile
xi362 net2303 net2501 net2504 net2498 net2497 net2503 net2502 net2304 vdd vss unit_coupling_tile
xi361 net2307 net2507 net2506 net2504 net2503 net2505 net2508 net2308 vdd vss unit_coupling_tile
xi360 net2311 net2511 net2510 net2506 net2505 net2509 net2512 net2312 vdd vss unit_coupling_tile
xi359 net2315 net2515 net2514 net2510 net2509 net2513 net2516 net2316 vdd vss unit_coupling_tile
xi358 net2320 net2519 net2518 net2514 net2513 net2517 net2520 net2317 vdd vss unit_coupling_tile
xi357 net2323 net2524 net2523 net2518 net2517 net2522 net2521 net2324 vdd vss unit_coupling_tile
xi356 net2325 net2527 net2526 net2523 net2522 net2525 net2528 net2326 vdd vss unit_coupling_tile
xi355 net2331 net2529 net2532 net2526 net2525 net2531 net2530 net2332 vdd vss unit_coupling_tile
xi354 net2335 net2535 net2534 net2532 net2531 net2533 net2536 net2336 vdd vss unit_coupling_tile
xi353 net2339 net2539 net2538 net2534 net2533 net2537 net2540 net2340 vdd vss unit_coupling_tile
xi352 net2343 net2543 net2542 net2538 net2537 net2541 net2544 net2344 vdd vss unit_coupling_tile
xi351 net2348 net2547 net2546 net2542 net2541 net2545 net2548 net2345 vdd vss unit_coupling_tile
xi350 net2351 net2552 net2551 net2546 net2545 net2550 net2549 net2352 vdd vss unit_coupling_tile
xi349 net2355 net2555 net2554 net96 net96 net2553 net2556 net2356 vdd vss unit_coupling_tile
xi348 net2357 net2559 net2558 net2554 net2553 net2557 net2560 net2358 vdd vss unit_coupling_tile
xi347 net2363 net2561 net2564 net2558 net2557 net2563 net2562 net2364 vdd vss unit_coupling_tile
xi346 net2367 net2567 net2566 net2564 net2563 net2565 net2568 net2368 vdd vss unit_coupling_tile
xi345 net2371 net2571 net2570 net2566 net2565 net2569 net2572 net2372 vdd vss unit_coupling_tile
xi344 net2376 net2575 net2574 net2570 net2569 net2573 net2576 net2373 vdd vss unit_coupling_tile
xi342 net2386 net2581 net2579 net2580 net2583 net2578 net2582 net2385 vdd vss unit_coupling_tile
xi341 net2382 net2587 net2586 net2579 net2578 net2585 net2588 net2383 vdd vss unit_coupling_tile
xi340 net2391 net2589 net2592 net2586 net2585 net2591 net2590 net2392 vdd vss unit_coupling_tile
xi339 net2395 net2595 net2594 net2592 net2591 net2593 net2596 net2396 vdd vss unit_coupling_tile
xi338 net2399 net2599 net2598 net2594 net2593 net2597 net2600 net2400 vdd vss unit_coupling_tile
xi337 net2404 net2603 net2602 net2598 net2597 net2601 net2604 net2401 vdd vss unit_coupling_tile
xi336 net2407 net2608 net2607 net2602 net2601 net2606 net2605 net2408 vdd vss unit_coupling_tile
xi335 net2411 net2611 net2610 net2607 net2606 net2609 net2612 net2412 vdd vss unit_coupling_tile
xi334 net2413 net2615 net2614 net2610 net2609 net2613 net2616 net2414 vdd vss unit_coupling_tile
xi333 net2419 net2617 net2620 net2614 net2613 net2619 net2618 net2420 vdd vss unit_coupling_tile
xi332 net2423 net2623 net2622 net2620 net2619 net2621 net2624 net2424 vdd vss unit_coupling_tile
xi331 net2427 net2627 net2626 net2622 net2621 net2625 net2628 net2428 vdd vss unit_coupling_tile
xi330 net2431 net2631 net2630 net2626 net2625 net2629 net2632 net2432 vdd vss unit_coupling_tile
xi329 net2436 net2635 net2634 net2630 net2629 net2633 net2636 net2433 vdd vss unit_coupling_tile
xi328 net2439 net2640 net2639 net2634 net2633 net2638 net2637 net2440 vdd vss unit_coupling_tile
xi327 net2441 net2643 net2642 net2639 net2638 net2641 net2644 net2442 vdd vss unit_coupling_tile
xi326 net2447 net2645 net2648 net2642 net2641 net2647 net2646 net2448 vdd vss unit_coupling_tile
xi325 net2451 net2651 net2650 net2648 net2647 net2649 net2652 net2452 vdd vss unit_coupling_tile
xi324 net2455 net2655 net2654 net2650 net2649 net2653 net2656 net2456 vdd vss unit_coupling_tile
xi323 net2459 net2659 net2658 net2654 net2653 net2657 net2660 net2460 vdd vss unit_coupling_tile
xi322 net2464 net2663 net2662 net2658 net2657 net2661 net2664 net2461 vdd vss unit_coupling_tile
xi321 net2467 net2668 net2667 net2662 net2661 net2666 net2665 net2468 vdd vss unit_coupling_tile
xi320 net2471 net2671 net2670 net2667 net2666 net2669 net2672 net2472 vdd vss unit_coupling_tile
xi319 net2473 net2675 net2674 net2670 net2669 net2673 net2676 net2474 vdd vss unit_coupling_tile
xi318 net2479 net2677 net2680 net2674 net2673 net2679 net2678 net2480 vdd vss unit_coupling_tile
xi317 net2483 net2683 net2682 net2680 net2679 net2681 net2684 net2484 vdd vss unit_coupling_tile
xi316 net2487 net2687 net2686 net2682 net2681 net2685 net2688 net2488 vdd vss unit_coupling_tile
xi315 net2492 net2691 net2690 net2686 net2685 net2689 net2692 net2489 vdd vss unit_coupling_tile
xi314 net2495 net2696 net2695 net2690 net2689 net2694 net2693 net2496 vdd vss unit_coupling_tile
xi313 net2499 net2699 net2698 net2695 net2694 net2697 net2700 net2500 vdd vss unit_coupling_tile
xi312 net2501 net2703 net2702 net2698 net2697 net2701 net2704 net2502 vdd vss unit_coupling_tile
xi311 net2507 net2705 net2708 net2702 net2701 net2707 net2706 net2508 vdd vss unit_coupling_tile
xi310 net2511 net2711 net2710 net2708 net2707 net2709 net2712 net2512 vdd vss unit_coupling_tile
xi309 net2515 net2715 net2714 net2710 net2709 net2713 net2716 net2516 vdd vss unit_coupling_tile
xi308 net2519 net2719 net2718 net2714 net2713 net2717 net2720 net2520 vdd vss unit_coupling_tile
xi307 net2524 net2723 net2722 net2718 net2717 net2721 net2724 net2521 vdd vss unit_coupling_tile
xi306 net2527 net2728 net2727 net2722 net2721 net2726 net2725 net2528 vdd vss unit_coupling_tile
xi305 net2529 net2731 net2730 net2727 net2726 net2729 net2732 net2530 vdd vss unit_coupling_tile
xi304 net2535 net2733 net2736 net2730 net2729 net2735 net2734 net2536 vdd vss unit_coupling_tile
xi303 net2539 net2739 net2738 net2736 net2735 net2737 net2740 net2540 vdd vss unit_coupling_tile
xi302 net2543 net2743 net2742 net2738 net2737 net2741 net2744 net2544 vdd vss unit_coupling_tile
xi301 net2547 net2747 net2746 net2742 net2741 net2745 net2748 net2548 vdd vss unit_coupling_tile
xi300 net2552 net2751 net2750 net2746 net2745 net2749 net2752 net2549 vdd vss unit_coupling_tile
xi299 net2555 net2756 net2755 net97 net97 net2754 net2753 net2556 vdd vss unit_coupling_tile
xi298 net2559 net2759 net2758 net2755 net2754 net2757 net2760 net2560 vdd vss unit_coupling_tile
xi297 net2561 net2763 net2762 net2758 net2757 net2761 net2764 net2562 vdd vss unit_coupling_tile
xi296 net2567 net2765 net2768 net2762 net2761 net2767 net2766 net2568 vdd vss unit_coupling_tile
xi295 net2571 net2771 net2770 net2768 net2767 net2769 net2772 net2572 vdd vss unit_coupling_tile
xi293 net2584 net2779 net2778 net2775 net2776 net2777 net2780 net2577 vdd vss unit_coupling_tile
xi292 net2581 net2784 net2783 net2778 net2777 net2782 net2781 net2582 vdd vss unit_coupling_tile
xi291 net2587 net2787 net2786 net2783 net2782 net2785 net2788 net2588 vdd vss unit_coupling_tile
xi290 net2589 net2791 net2790 net2786 net2785 net2789 net2792 net2590 vdd vss unit_coupling_tile
xi289 net2595 net2793 net2796 net2790 net2789 net2795 net2794 net2596 vdd vss unit_coupling_tile
xi288 net2599 net2799 net2798 net2796 net2795 net2797 net2800 net2600 vdd vss unit_coupling_tile
xi287 net2603 net2803 net2802 net2798 net2797 net2801 net2804 net2604 vdd vss unit_coupling_tile
xi286 net2608 net2807 net2806 net2802 net2801 net2805 net2808 net2605 vdd vss unit_coupling_tile
xi285 net2611 net2812 net2811 net2806 net2805 net2810 net2809 net2612 vdd vss unit_coupling_tile
xi284 net2615 net2815 net2814 net2811 net2810 net2813 net2816 net2616 vdd vss unit_coupling_tile
xi283 net2617 net2819 net2818 net2814 net2813 net2817 net2820 net2618 vdd vss unit_coupling_tile
xi282 net2623 net2821 net2824 net2818 net2817 net2823 net2822 net2624 vdd vss unit_coupling_tile
xi281 net2627 net2827 net2826 net2824 net2823 net2825 net2828 net2628 vdd vss unit_coupling_tile
xi280 net2631 net2831 net2830 net2826 net2825 net2829 net2832 net2632 vdd vss unit_coupling_tile
xi279 net2635 net2835 net2834 net2830 net2829 net2833 net2836 net2636 vdd vss unit_coupling_tile
xi278 net2640 net2840 net2841 net2834 net2833 net2837 net2839 net2637 vdd vss unit_coupling_tile
xi277 net2643 net2848 net2845 net2841 net2837 net2842 net2838 net2644 vdd vss unit_coupling_tile
xi276 net2645 net2844 net2846 net2845 net2842 net2847 net2843 net2646 vdd vss unit_coupling_tile
xi275 net2651 net2850 net2855 net2846 net2847 net2852 net2849 net2652 vdd vss unit_coupling_tile
xi274 net2655 net2854 net2856 net2855 net2852 net2851 net2853 net2656 vdd vss unit_coupling_tile
xi273 net2659 net2864 net2860 net2856 net2851 net2857 net2863 net2660 vdd vss unit_coupling_tile
xi272 net2663 net2859 net2861 net2860 net2857 net2862 net2858 net2664 vdd vss unit_coupling_tile
xi271 net2668 net2868 net2869 net2861 net2862 net2865 net2867 net2665 vdd vss unit_coupling_tile
xi270 net2671 net2876 net2873 net2869 net2865 net2870 net2866 net2672 vdd vss unit_coupling_tile
xi269 net2675 net2872 net2874 net2873 net2870 net2875 net2871 net2676 vdd vss unit_coupling_tile
xi268 net2677 net2882 net2880 net2874 net2875 net2877 net2881 net2678 vdd vss unit_coupling_tile
xi267 net2683 net2879 net2887 net2880 net2877 net2884 net2878 net2684 vdd vss unit_coupling_tile
xi266 net2687 net2886 net2888 net2887 net2884 net2883 net2885 net2688 vdd vss unit_coupling_tile
xi265 net2691 net2890 net2891 net2888 net2883 net2892 net2889 net2692 vdd vss unit_coupling_tile
xi264 net2696 net2896 net2897 net2891 net2892 net2893 net2895 net2693 vdd vss unit_coupling_tile
xi263 net2699 net2904 net2901 net2897 net2893 net2898 net2894 net2700 vdd vss unit_coupling_tile
xi262 net2703 net2900 net2902 net2901 net2898 net2903 net2899 net2704 vdd vss unit_coupling_tile
xi261 net2705 net2910 net2908 net2902 net2903 net2905 net2909 net2706 vdd vss unit_coupling_tile
xi260 net2711 net2907 net2915 net2908 net2905 net2912 net2906 net2712 vdd vss unit_coupling_tile
xi259 net2715 net2914 net2916 net2915 net2912 net2911 net2913 net2716 vdd vss unit_coupling_tile
xi258 net2719 net2924 net2920 net2916 net2911 net2917 net2923 net2720 vdd vss unit_coupling_tile
xi257 net2723 net2919 net2921 net2920 net2917 net2922 net2918 net2724 vdd vss unit_coupling_tile
xi256 net2728 net2928 net2929 net2921 net2922 net2925 net2927 net2725 vdd vss unit_coupling_tile
xi255 net2731 net2930 net2931 net2929 net2925 net2932 net2926 net2732 vdd vss unit_coupling_tile
xi254 net2733 net2938 net2936 net2931 net2932 net2933 net2937 net2734 vdd vss unit_coupling_tile
xi253 net2739 net2935 net2943 net2936 net2933 net2940 net2934 net2740 vdd vss unit_coupling_tile
xi252 net2743 net2942 net2944 net2943 net2940 net2939 net2941 net2744 vdd vss unit_coupling_tile
xi251 net2747 net2952 net2948 net2944 net2939 net2945 net2951 net2748 vdd vss unit_coupling_tile
xi250 net2751 net2947 net2949 net2948 net2945 net2950 net2946 net2752 vdd vss unit_coupling_tile
xi249 net2756 net2956 net2957 net98 net98 net2953 net2955 net2753 vdd vss unit_coupling_tile
xi248 net2759 net2964 net2961 net2957 net2953 net2958 net2954 net2760 vdd vss unit_coupling_tile
xi247 net2763 net2960 net2962 net2961 net2958 net2963 net2959 net2764 vdd vss unit_coupling_tile
xi246 net2765 net2966 net2967 net2962 net2963 net2968 net2965 net2766 vdd vss unit_coupling_tile
xi244 net2774 net2979 net2975 net2972 net2971 net2973 net2978 net2773 vdd vss unit_coupling_tile
xi243 net2779 net378 net2976 net2975 net2973 net2977 net2974 net2780 vdd vss unit_coupling_tile
xi242 net2784 net372 net2981 net2976 net2977 net2980 net371 net2781 vdd vss unit_coupling_tile
xi241 net2787 net389 net2983 net2981 net2980 net2982 net388 net2788 vdd vss unit_coupling_tile
xi240 net2791 net386 net2984 net2983 net2982 net2985 net385 net2792 vdd vss unit_coupling_tile
xi239 net2793 net397 net2987 net2984 net2985 net2986 net396 net2794 vdd vss unit_coupling_tile
xi238 net2799 net413 net2990 net2987 net2986 net2989 net412 net2800 vdd vss unit_coupling_tile
xi237 net2803 net408 net2991 net2990 net2989 net2988 net407 net2804 vdd vss unit_coupling_tile
xi236 net2807 net420 net2993 net2991 net2988 net2992 net419 net2808 vdd vss unit_coupling_tile
xi235 net2812 net435 net2994 net2993 net2992 net2995 net417 net2809 vdd vss unit_coupling_tile
xi234 net2815 net429 net2997 net2994 net2995 net2996 net428 net2816 vdd vss unit_coupling_tile
xi233 net2819 net439 net2998 net2997 net2996 net2999 net438 net2820 vdd vss unit_coupling_tile
xi232 net2821 net507 net3001 net2998 net2999 net3000 net506 net2822 vdd vss unit_coupling_tile
xi231 net2827 net523 net3004 net3001 net3000 net3003 net522 net2828 vdd vss unit_coupling_tile
xi230 net2831 net518 net3005 net3004 net3003 net3002 net517 net2832 vdd vss unit_coupling_tile
xi229 net2835 net530 net3007 net3005 net3002 net3006 net529 net2836 vdd vss unit_coupling_tile
xi228 net2840 net545 net3008 net3007 net3006 net3009 net527 net2839 vdd vss unit_coupling_tile
xi227 net2848 net539 net3011 net3008 net3009 net3010 net538 net2838 vdd vss unit_coupling_tile
xi226 net2844 net553 net3013 net3011 net3010 net3012 net552 net2843 vdd vss unit_coupling_tile
xi225 net2850 net550 net3014 net3013 net3012 net3015 net549 net2849 vdd vss unit_coupling_tile
xi224 net2854 net561 net3018 net3014 net3015 net3017 net560 net2853 vdd vss unit_coupling_tile
xi223 net2864 net571 net3019 net3018 net3017 net3016 net570 net2863 vdd vss unit_coupling_tile
xi222 net2859 net809 net3021 net3019 net3016 net3020 net808 net2858 vdd vss unit_coupling_tile
xi221 net2868 net822 net3022 net3021 net3020 net3023 net806 net2867 vdd vss unit_coupling_tile
xi220 net2876 net816 net3025 net3022 net3023 net3024 net815 net2866 vdd vss unit_coupling_tile
xi219 net2872 net830 net3027 net3025 net3024 net3026 net829 net2871 vdd vss unit_coupling_tile
xi218 net2882 net827 net3028 net3027 net3026 net3029 net826 net2881 vdd vss unit_coupling_tile
xi217 net2879 net838 net3031 net3028 net3029 net3030 net837 net2878 vdd vss unit_coupling_tile
xi216 net2886 net854 net3034 net3031 net3030 net3033 net853 net2885 vdd vss unit_coupling_tile
xi215 net2890 net849 net3035 net3034 net3033 net3032 net848 net2889 vdd vss unit_coupling_tile
xi214 net2896 net861 net3036 net3035 net3032 net3037 net860 net2895 vdd vss unit_coupling_tile
xi213 net2904 net866 net3039 net3036 net3037 net3038 net858 net2894 vdd vss unit_coupling_tile
xi212 net2900 net768 net3041 net3039 net3038 net3040 net767 net2899 vdd vss unit_coupling_tile
xi211 net2910 net765 net3042 net3041 net3040 net3043 net764 net2909 vdd vss unit_coupling_tile
xi210 net2907 net775 net3045 net3042 net3043 net3044 net774 net2906 vdd vss unit_coupling_tile
xi209 net2914 net784 net3048 net3045 net3044 net3047 net783 net2913 vdd vss unit_coupling_tile
xi208 net2924 net781 net3049 net3048 net3047 net3046 net780 net2923 vdd vss unit_coupling_tile
xi207 net2919 net789 net3051 net3049 net3046 net3050 net788 net2918 vdd vss unit_coupling_tile
xi206 net2928 net798 net3052 net3051 net3050 net3053 net786 net2927 vdd vss unit_coupling_tile
xi205 net2930 net794 net3055 net3052 net3053 net3054 net793 net2926 vdd vss unit_coupling_tile
xi204 net2938 net803 net3056 net3055 net3054 net3057 net802 net2937 vdd vss unit_coupling_tile
xi203 net2935 net801 net3059 net3056 net3057 net3058 net800 net2934 vdd vss unit_coupling_tile
xi202 net2942 net692 net3062 net3059 net3058 net3061 net691 net2941 vdd vss unit_coupling_tile
xi201 net2952 net688 net3063 net3062 net3061 net3060 net687 net2951 vdd vss unit_coupling_tile
xi200 net2947 net697 net3066 net3063 net3060 net3067 net696 net2946 vdd vss unit_coupling_tile
xi199 net2956 net707 net3064 net99 net99 net3065 net694 net2955 vdd vss unit_coupling_tile
xi198 net2964 net703 net3069 net3064 net3065 net3068 net702 net2954 vdd vss unit_coupling_tile
xi197 net2960 net712 net3070 net3069 net3068 net3071 net711 net2959 vdd vss unit_coupling_tile
xi195 net2970 net716 net3075 net3072 net3073 net3074 net715 net2969 vdd vss unit_coupling_tile
xi194 net2979 net723 net381 net3075 net3074 net3076 net722 net2978 vdd vss unit_coupling_tile
xi193 net378 net380 net375 net381 net3076 net370 net379 net2974 vdd vss unit_coupling_tile
xi192 net372 net374 net376 net375 net370 net377 net373 net371 vdd vss unit_coupling_tile
xi191 net389 net391 net392 net376 net377 net384 net390 net388 vdd vss unit_coupling_tile
xi190 net386 net405 net400 net392 net384 net395 net387 net385 vdd vss unit_coupling_tile
xi189 net397 net399 net401 net400 net395 net402 net398 net396 vdd vss unit_coupling_tile
xi188 net413 net415 net411 net401 net402 net406 net414 net412 vdd vss unit_coupling_tile
xi187 net408 net410 net423 net411 net406 net418 net409 net407 vdd vss unit_coupling_tile
xi186 net420 net422 net424 net423 net418 net416 net421 net419 vdd vss unit_coupling_tile
xi185 net435 net437 net432 net424 net416 net427 net436 net417 vdd vss unit_coupling_tile
xi184 net429 net431 net433 net432 net427 net434 net430 net428 vdd vss unit_coupling_tile
xi183 net439 net515 net510 net433 net434 net505 net440 net438 vdd vss unit_coupling_tile
xi182 net507 net509 net511 net510 net505 net512 net508 net506 vdd vss unit_coupling_tile
xi181 net523 net525 net521 net511 net512 net516 net524 net522 vdd vss unit_coupling_tile
xi180 net518 net520 net533 net521 net516 net528 net519 net517 vdd vss unit_coupling_tile
xi179 net530 net532 net534 net533 net528 net526 net531 net529 vdd vss unit_coupling_tile
xi178 net545 net547 net542 net534 net526 net537 net546 net527 vdd vss unit_coupling_tile
xi177 net539 net541 net543 net542 net537 net544 net540 net538 vdd vss unit_coupling_tile
xi176 net553 net555 net556 net543 net544 net548 net554 net552 vdd vss unit_coupling_tile
xi175 net550 net569 net564 net556 net548 net559 net551 net549 vdd vss unit_coupling_tile
xi174 net561 net563 net565 net564 net559 net566 net562 net560 vdd vss unit_coupling_tile
xi173 net571 net573 net810 net565 net566 net807 net572 net570 vdd vss unit_coupling_tile
xi172 net809 net683 net811 net810 net807 net805 net682 net808 vdd vss unit_coupling_tile
xi171 net822 net824 net819 net811 net805 net814 net823 net806 vdd vss unit_coupling_tile
xi170 net816 net818 net820 net819 net814 net821 net817 net815 vdd vss unit_coupling_tile
xi169 net830 net832 net833 net820 net821 net825 net831 net829 vdd vss unit_coupling_tile
xi168 net827 net846 net841 net833 net825 net836 net828 net826 vdd vss unit_coupling_tile
xi167 net838 net840 net842 net841 net836 net843 net839 net837 vdd vss unit_coupling_tile
xi166 net854 net856 net852 net842 net843 net847 net855 net853 vdd vss unit_coupling_tile
xi165 net849 net851 net864 net852 net847 net859 net850 net848 vdd vss unit_coupling_tile
xi164 net861 net863 net865 net864 net859 net857 net862 net860 vdd vss unit_coupling_tile
xi163 net866 net868 net771 net865 net857 net766 net867 net858 vdd vss unit_coupling_tile
xi162 net768 net770 net772 net771 net766 net763 net769 net767 vdd vss unit_coupling_tile
xi161 net765 net580 net776 net772 net763 net773 net579 net764 vdd vss unit_coupling_tile
xi160 net775 net576 net777 net776 net773 net778 net575 net774 vdd vss unit_coupling_tile
xi159 net784 net589 net782 net777 net778 net779 net588 net783 vdd vss unit_coupling_tile
xi158 net781 net605 net790 net782 net779 net787 net604 net780 vdd vss unit_coupling_tile
xi157 net789 net600 net791 net790 net787 net785 net599 net788 vdd vss unit_coupling_tile
xi156 net798 net612 net795 net791 net785 net792 net611 net786 vdd vss unit_coupling_tile
xi155 net794 net627 net796 net795 net792 net797 net609 net793 vdd vss unit_coupling_tile
xi154 net803 net621 net804 net796 net797 net799 net620 net802 vdd vss unit_coupling_tile
xi153 net801 net635 net693 net804 net799 net690 net634 net800 vdd vss unit_coupling_tile
xi152 net692 net632 net689 net693 net690 net686 net631 net691 vdd vss unit_coupling_tile
xi151 net688 net309 net698 net689 net686 net695 net308 net687 vdd vss unit_coupling_tile
xi150 net697 net303 net699 net698 net695 net700 net302 net696 vdd vss unit_coupling_tile
xi149 net707 net316 net704 net100 net100 net701 net315 net694 vdd vss unit_coupling_tile
xi148 net703 net332 net705 net704 net701 net706 net323 net702 vdd vss unit_coupling_tile
xi146 net710 net340 net717 net713 net708 net714 net339 net709 vdd vss unit_coupling_tile
xi145 net716 net337 net718 net717 net714 net719 net336 net715 vdd vss unit_coupling_tile
xi144 net723 net348 net721 net718 net719 net720 net347 net722 vdd vss unit_coupling_tile
xi143 net380 net364 net725 net721 net720 net724 net363 net379 vdd vss unit_coupling_tile
xi142 net374 net359 net728 net725 net724 net726 net358 net373 vdd vss unit_coupling_tile
xi141 net391 net727 net729 net728 net726 net730 net368 net390 vdd vss unit_coupling_tile
xi140 net405 net734 net735 net729 net730 net731 net733 net387 vdd vss unit_coupling_tile
xi139 net399 net742 net739 net735 net731 net736 net732 net398 vdd vss unit_coupling_tile
xi138 net415 net738 net740 net739 net736 net741 net737 net414 vdd vss unit_coupling_tile
xi137 net410 net748 net746 net740 net741 net743 net747 net409 vdd vss unit_coupling_tile
xi136 net422 net745 net753 net746 net743 net750 net744 net421 vdd vss unit_coupling_tile
xi135 net437 net752 net754 net753 net750 net749 net751 net436 vdd vss unit_coupling_tile
xi134 net431 net761 net758 net754 net749 net755 net760 net430 vdd vss unit_coupling_tile
xi133 net515 net757 net647 net758 net755 net759 net756 net440 vdd vss unit_coupling_tile
xi132 net509 net646 net643 net647 net759 net640 net762 net508 vdd vss unit_coupling_tile
xi131 net525 net642 net644 net643 net640 net645 net641 net524 vdd vss unit_coupling_tile
xi130 net520 net653 net651 net644 net645 net648 net652 net519 vdd vss unit_coupling_tile
xi129 net532 net650 net658 net651 net648 net655 net649 net531 vdd vss unit_coupling_tile
xi128 net547 net657 net659 net658 net655 net654 net656 net546 vdd vss unit_coupling_tile
xi127 net541 net667 net663 net659 net654 net660 net666 net540 vdd vss unit_coupling_tile
xi126 net555 net662 net664 net663 net660 net665 net661 net554 vdd vss unit_coupling_tile
xi125 net569 net671 net672 net664 net665 net668 net670 net551 vdd vss unit_coupling_tile
xi124 net563 net681 net676 net672 net668 net673 net669 net562 vdd vss unit_coupling_tile
xi123 net573 net675 net677 net676 net673 net678 net674 net572 vdd vss unit_coupling_tile
xi122 net683 net685 net873 net677 net678 net870 net684 net682 vdd vss unit_coupling_tile
xi121 net824 net872 net874 net873 net870 net869 net871 net823 vdd vss unit_coupling_tile
xi120 net818 net882 net878 net874 net869 net875 net881 net817 vdd vss unit_coupling_tile
xi119 net832 net877 net879 net878 net875 net880 net876 net831 vdd vss unit_coupling_tile
xi118 net846 net886 net887 net879 net880 net883 net885 net828 vdd vss unit_coupling_tile
xi117 net840 net894 net891 net887 net883 net888 net884 net839 vdd vss unit_coupling_tile
xi116 net856 net890 net892 net891 net888 net893 net889 net855 vdd vss unit_coupling_tile
xi115 net851 net900 net898 net892 net893 net895 net899 net850 vdd vss unit_coupling_tile
xi114 net863 net897 net905 net898 net895 net902 net896 net862 vdd vss unit_coupling_tile
xi113 net868 net904 net906 net905 net902 net901 net903 net867 vdd vss unit_coupling_tile
xi112 net770 net908 net583 net906 net901 net578 net907 net769 vdd vss unit_coupling_tile
xi111 net580 net582 net584 net583 net578 net574 net581 net579 vdd vss unit_coupling_tile
xi110 net576 net597 net592 net584 net574 net587 net577 net575 vdd vss unit_coupling_tile
xi109 net589 net591 net593 net592 net587 net594 net590 net588 vdd vss unit_coupling_tile
xi108 net605 net607 net603 net593 net594 net598 net606 net604 vdd vss unit_coupling_tile
xi107 net600 net602 net615 net603 net598 net610 net601 net599 vdd vss unit_coupling_tile
xi106 net612 net614 net616 net615 net610 net608 net613 net611 vdd vss unit_coupling_tile
xi105 net627 net629 net624 net616 net608 net619 net628 net609 vdd vss unit_coupling_tile
xi104 net621 net623 net625 net624 net619 net626 net622 net620 vdd vss unit_coupling_tile
xi103 net635 net637 net638 net625 net626 net630 net636 net634 vdd vss unit_coupling_tile
xi102 net632 net639 net312 net638 net630 net307 net633 net631 vdd vss unit_coupling_tile
xi101 net309 net311 net306 net312 net307 net301 net310 net308 vdd vss unit_coupling_tile
xi100 net303 net305 net321 net306 net301 net322 net304 net302 vdd vss unit_coupling_tile
xi99 net316 net318 net319 net101 net101 net320 net317 net315 vdd vss unit_coupling_tile
xi97 net326 net328 net330 net329 net324 net331 net327 net325 vdd vss unit_coupling_tile
xi96 net340 net342 net343 net330 net331 net335 net341 net339 vdd vss unit_coupling_tile
xi95 net337 net356 net351 net343 net335 net346 net338 net336 vdd vss unit_coupling_tile
xi94 net348 net350 net352 net351 net346 net353 net349 net347 vdd vss unit_coupling_tile
xi93 net364 net366 net362 net352 net353 net357 net365 net363 vdd vss unit_coupling_tile
xi92 net359 net361 net369 net362 net357 net367 net360 net358 vdd vss unit_coupling_tile
xi91 net727 net1361 net1775 net369 net367 net1773 net1362 net368 vdd vss unit_coupling_tile
xi90 net734 net1774 net1776 net1775 net1773 net1777 net1365 net733 vdd vss unit_coupling_tile
xi89 net742 net1781 net1782 net1776 net1777 net1778 net1780 net732 vdd vss unit_coupling_tile
xi88 net738 net1789 net1786 net1782 net1778 net1783 net1779 net737 vdd vss unit_coupling_tile
xi87 net748 net1785 net1787 net1786 net1783 net1788 net1784 net747 vdd vss unit_coupling_tile
xi86 net745 net1795 net1793 net1787 net1788 net1790 net1794 net744 vdd vss unit_coupling_tile
xi85 net752 net1792 net1800 net1793 net1790 net1797 net1791 net751 vdd vss unit_coupling_tile
xi84 net761 net1799 net1801 net1800 net1797 net1796 net1798 net760 vdd vss unit_coupling_tile
xi83 net757 net1809 net1805 net1801 net1796 net1802 net1808 net756 vdd vss unit_coupling_tile
xi82 net646 net1804 net1806 net1805 net1802 net1807 net1803 net762 vdd vss unit_coupling_tile
xi81 net642 net1817 net1814 net1806 net1807 net1811 net1810 net641 vdd vss unit_coupling_tile
xi80 net653 net1813 net1815 net1814 net1811 net1816 net1812 net652 vdd vss unit_coupling_tile
xi79 net650 net1145 net1819 net1815 net1816 net1818 net1146 net649 vdd vss unit_coupling_tile
xi78 net657 net1149 net1822 net1819 net1818 net1821 net1150 net656 vdd vss unit_coupling_tile
xi77 net667 net1151 net1823 net1822 net1821 net1820 net1152 net666 vdd vss unit_coupling_tile
xi76 net662 net1157 net1825 net1823 net1820 net1824 net1158 net661 vdd vss unit_coupling_tile
xi75 net671 net1162 net1826 net1825 net1824 net1827 net1159 net670 vdd vss unit_coupling_tile
xi74 net681 net1165 net1829 net1826 net1827 net1828 net1166 net669 vdd vss unit_coupling_tile
xi73 net675 net1169 net1831 net1829 net1828 net1830 net1170 net674 vdd vss unit_coupling_tile
xi72 net685 net1171 net1832 net1831 net1830 net1833 net1172 net684 vdd vss unit_coupling_tile
xi71 net872 net1177 net913 net1832 net1833 net910 net1178 net871 vdd vss unit_coupling_tile
xi70 net882 net912 net914 net913 net910 net909 net911 net881 vdd vss unit_coupling_tile
xi69 net877 net917 net916 net914 net909 net915 net918 net876 vdd vss unit_coupling_tile
xi68 net886 net921 net920 net916 net915 net919 net922 net885 vdd vss unit_coupling_tile
xi67 net894 net925 net924 net920 net919 net923 net926 net884 vdd vss unit_coupling_tile
xi66 net890 net930 net929 net924 net923 net928 net927 net889 vdd vss unit_coupling_tile
xi65 net900 net933 net932 net929 net928 net931 net934 net899 vdd vss unit_coupling_tile
xi64 net897 net937 net936 net932 net931 net935 net938 net896 vdd vss unit_coupling_tile
xi63 net904 net939 net942 net936 net935 net941 net940 net903 vdd vss unit_coupling_tile
xi62 net908 net945 net944 net942 net941 net943 net946 net907 vdd vss unit_coupling_tile
xi61 net582 net949 net948 net944 net943 net947 net950 net581 vdd vss unit_coupling_tile
xi60 net597 net972 net976 net948 net947 net975 net968 net577 vdd vss unit_coupling_tile
xi59 net591 net980 net979 net976 net975 net978 net977 net590 vdd vss unit_coupling_tile
xi58 net607 net983 net982 net979 net978 net981 net984 net606 vdd vss unit_coupling_tile
xi57 net602 net987 net986 net982 net981 net985 net988 net601 vdd vss unit_coupling_tile
xi56 net614 net989 net992 net986 net985 net991 net990 net613 vdd vss unit_coupling_tile
xi55 net629 net995 net994 net992 net991 net993 net996 net628 vdd vss unit_coupling_tile
xi54 net623 net999 net998 net994 net993 net997 net1000 net622 vdd vss unit_coupling_tile
xi53 net637 net1003 net1002 net998 net997 net1001 net1004 net636 vdd vss unit_coupling_tile
xi52 net639 net1007 net1006 net1002 net1001 net1005 net1008 net633 vdd vss unit_coupling_tile
xi51 net311 net1012 net1011 net1006 net1005 net1010 net1009 net310 vdd vss unit_coupling_tile
xi50 net305 net1255 net1344 net1011 net1010 net1343 net1254 net304 vdd vss unit_coupling_tile
xi48 net334 net51 net1346 net1347 net1348 net1345 net51 net333 vdd vss unit_coupling_tile
xi47 net328 net50 net1350 net1346 net1345 net1349 net50 net327 vdd vss unit_coupling_tile
xi46 net342 net49 net1352 net1350 net1349 net1351 net49 net341 vdd vss unit_coupling_tile
xi45 net356 net48 net1354 net1352 net1351 net1353 net48 net338 vdd vss unit_coupling_tile
xi44 net350 net47 net1356 net1354 net1353 net1355 net47 net349 vdd vss unit_coupling_tile
xi43 net366 net46 net1358 net1356 net1355 net1357 net46 net365 vdd vss unit_coupling_tile
xi42 net361 net45 net1360 net1358 net1357 net1359 net45 net360 vdd vss unit_coupling_tile
xi41 net1361 net44 net1364 net1360 net1359 net1363 net44 net1362 vdd vss unit_coupling_tile
xi40 net1774 net43 net1895 net1364 net1363 net1894 net43 net1365 vdd vss unit_coupling_tile
xi39 net1781 net42 net1897 net1895 net1894 net1896 net42 net1780 vdd vss unit_coupling_tile
xi38 net1789 net41 net1899 net1897 net1896 net1898 net41 net1779 vdd vss unit_coupling_tile
xi37 net1785 net40 net1901 net1899 net1898 net1900 net40 net1784 vdd vss unit_coupling_tile
xi36 net1795 net39 net1903 net1901 net1900 net1902 net39 net1794 vdd vss unit_coupling_tile
xi35 net1792 net38 net1905 net1903 net1902 net1904 net38 net1791 vdd vss unit_coupling_tile
xi34 net1799 net37 net1907 net1905 net1904 net1906 net37 net1798 vdd vss unit_coupling_tile
xi33 net1809 net36 net1909 net1907 net1906 net1908 net36 net1808 vdd vss unit_coupling_tile
xi32 net1804 net35 net1911 net1909 net1908 net1910 net35 net1803 vdd vss unit_coupling_tile
xi31 net1817 net34 net1142 net1911 net1910 net1912 net34 net1810 vdd vss unit_coupling_tile
xi30 net1813 net33 net1141 net1142 net1912 net1140 net33 net1812 vdd vss unit_coupling_tile
xi29 net1145 net32 net1144 net1141 net1140 net1143 net32 net1146 vdd vss unit_coupling_tile
xi28 net1149 net31 net1148 net1144 net1143 net1147 net31 net1150 vdd vss unit_coupling_tile
xi27 net1151 net30 net1154 net1148 net1147 net1153 net30 net1152 vdd vss unit_coupling_tile
xi26 net1157 net29 net1156 net1154 net1153 net1155 net29 net1158 vdd vss unit_coupling_tile
xi25 net1162 net28 net1161 net1156 net1155 net1160 net28 net1159 vdd vss unit_coupling_tile
xi24 net1165 net27 net1164 net1161 net1160 net1163 net27 net1166 vdd vss unit_coupling_tile
xi23 net1169 net26 net1168 net1164 net1163 net1167 net26 net1170 vdd vss unit_coupling_tile
xi22 net1171 net25 net1174 net1168 net1167 net1173 net25 net1172 vdd vss unit_coupling_tile
xi21 net1177 net24 net1176 net1174 net1173 net1175 net24 net1178 vdd vss unit_coupling_tile
xi20 net912 net23 net952 net1176 net1175 net951 net23 net911 vdd vss unit_coupling_tile
xi19 net917 net22 net954 net952 net951 net953 net22 net918 vdd vss unit_coupling_tile
xi18 net921 net21 net956 net954 net953 net955 net21 net922 vdd vss unit_coupling_tile
xi17 net925 net20 net958 net956 net955 net957 net20 net926 vdd vss unit_coupling_tile
xi16 net930 net19 net960 net958 net957 net959 net19 net927 vdd vss unit_coupling_tile
xi15 net933 net18 net962 net960 net959 net961 net18 net934 vdd vss unit_coupling_tile
xi14 net937 net17 net963 net962 net961 net964 net17 net938 vdd vss unit_coupling_tile
xi13 net939 net16 net966 net963 net964 net965 net16 net940 vdd vss unit_coupling_tile
xi12 net945 net15 net970 net966 net965 net969 net15 net946 vdd vss unit_coupling_tile
xi11 net949 net14 net971 net970 net969 net967 net14 net950 vdd vss unit_coupling_tile
xi10 net972 net13 net973 net971 net967 net974 net13 net968 vdd vss unit_coupling_tile
xi9 net980 net12 net1238 net973 net974 net1237 net12 net977 vdd vss unit_coupling_tile
xi8 net983 net11 net1240 net1238 net1237 net1239 net11 net984 vdd vss unit_coupling_tile
xi7 net987 net10 net1241 net1240 net1239 net1242 net10 net988 vdd vss unit_coupling_tile
xi6 net989 net9 net1244 net1241 net1242 net1243 net9 net990 vdd vss unit_coupling_tile
xi5 net995 net8 net1247 net1244 net1243 net1246 net8 net996 vdd vss unit_coupling_tile
xi4 net999 net7 net1248 net1247 net1246 net1245 net7 net1000 vdd vss unit_coupling_tile
xi3 net1003 net6 net1250 net1248 net1245 net1249 net6 net1004 vdd vss unit_coupling_tile
xi2 net1007 net5 net1251 net1250 net1249 net1252 net5 net1008 vdd vss unit_coupling_tile
xi1 net1012 net4 net1256 net1251 net1252 net1253 net4 net1009 vdd vss unit_coupling_tile
xi0 net1255 net3 net1257 net1256 net1253 net1258 net3 net1254 vdd vss unit_coupling_tile
xi2450 net10168 net9964 net10169 net10165 net10166 net10170 net9954 net10167 vdd vss short_tile
xi49 net318 net52 net1347 net102 net102 net1348 net52 net317 vdd vss short_tile
xi98 net332 net334 net329 net319 net320 net324 net333 net323 vdd vss short_tile
xi147 net712 net326 net713 net705 net706 net708 net325 net711 vdd vss short_tile
xi196 net2966 net710 net3072 net3070 net3071 net3073 net709 net2965 vdd vss short_tile
xi245 net2771 net2970 net2972 net2967 net2968 net2971 net2969 net2772 vdd vss short_tile
xi294 net2575 net2774 net2775 net2770 net2769 net2776 net2773 net2576 vdd vss short_tile
xi343 net2379 net2584 net2580 net2574 net2573 net2583 net2577 net2380 vdd vss short_tile
xi392 net2181 net2386 net2381 net2378 net2377 net2384 net2385 net2182 vdd vss short_tile
xi441 net1987 net2187 net2188 net2184 net2183 net2185 net2186 net1988 vdd vss short_tile
xi490 net1714 net1990 net1991 net1986 net1985 net1992 net1989 net1709 vdd vss short_tile
xi539 net1716 net1718 net1719 net1713 net1712 net1720 net1717 net1715 vdd vss short_tile
xi588 net1427 net1725 net1862 net1859 net1858 net1863 net1726 net1428 vdd vss short_tile
xi637 net1440 net1442 net1434 net1426 net1425 net1439 net1441 net1431 vdd vss short_tile
xi686 net3108 net1437 net3109 net3101 net3100 net3106 net1438 net3107 vdd vss short_tile
xi735 net3317 net3104 net3318 net3315 net3314 net3319 net3105 net3316 vdd vss short_tile
xi784 net3450 net3320 net3451 net3446 net3445 net3448 net3321 net3449 vdd vss short_tile
xi833 net3660 net3454 net3661 net3657 net3656 net3662 net3447 net3659 vdd vss short_tile
xi882 net3872 net3665 net3875 net3868 net3867 net3878 net3666 net3871 vdd vss short_tile
xi931 net4088 net3876 net4083 net4080 net4079 net4086 net3877 net4087 vdd vss short_tile
xi980 net4298 net4084 net4299 net4294 net4293 net4296 net4085 net4297 vdd vss short_tile
xi1029 net4430 net4300 net4432 net4431 net4428 net4427 net4295 net4429 vdd vss short_tile
xi1078 net4640 net4425 net4641 net4638 net4637 net4642 net4426 net4639 vdd vss short_tile
xi1127 net4852 net4645 net4858 net4849 net4850 net4855 net4646 net4851 vdd vss short_tile
xi1176 net5070 net4857 net5067 net5061 net5062 net5064 net4856 net5063 vdd vss short_tile
xi1225 net5279 net5066 net5280 net5272 net5273 net5275 net5065 net5278 vdd vss short_tile
xi1274 net5409 net5277 net5406 net5410 net5407 net5403 net5276 net5408 vdd vss short_tile
xi1323 net5620 net5405 net5621 net5617 net5618 net5615 net5404 net5619 vdd vss short_tile
xi1372 net5830 net5628 net5831 net5827 net5828 net5832 net5616 net5829 vdd vss short_tile
xi1421 net6042 net5837 net6046 net6039 net6040 net6043 net5836 net6041 vdd vss short_tile
xi1470 net6258 net6045 net6256 net6251 net6252 net6253 net6044 net6257 vdd vss short_tile
xi1519 net6388 net6255 net6385 net6389 net6463 net6382 net6254 net6464 vdd vss short_tile
xi1568 net6598 net6384 net6599 net6590 net6591 net6594 net6383 net6597 vdd vss short_tile
xi1617 net6807 net6596 net6808 net6804 net6805 net6809 net6595 net6806 vdd vss short_tile
xi1666 net7019 net6815 net7025 net7016 net7017 net7022 net6814 net7018 vdd vss short_tile
xi1715 net7236 net7024 net7234 net7228 net7229 net7231 net7023 net7230 vdd vss short_tile
xi1764 net7442 net7233 net7364 net7367 net7439 net7361 net7232 net7441 vdd vss short_tile
xi1813 net7577 net7363 net7575 net7569 net7570 net7572 net7362 net7576 vdd vss short_tile
xi1862 net7787 net7574 net7788 net7784 net7785 net7782 net7573 net7786 vdd vss short_tile
xi1911 net7997 net7795 net7998 net7994 net7995 net7999 net7783 net7996 vdd vss short_tile
xi1960 net8209 net8004 net8213 net8206 net8207 net8210 net8003 net8208 vdd vss short_tile
xi2009 net8421 net8212 net8346 net8418 net8419 net8343 net8211 net8420 vdd vss short_tile
xi2058 net8556 net8345 net8553 net8547 net8548 net8550 net8344 net8549 vdd vss short_tile
xi2107 net8767 net8552 net8768 net8760 net8761 net8763 net8551 net8766 vdd vss short_tile
xi2156 net8976 net8765 net8977 net8973 net8974 net8978 net8764 net8975 vdd vss short_tile
xi2205 net9188 net8984 net9194 net9185 net9186 net9191 net8983 net9187 vdd vss short_tile
xi2254 net9400 net9193 net9327 net9397 net9398 net9324 net9192 net9399 vdd vss short_tile
xi2303 net9532 net9326 net9536 net9529 net9530 net9533 net9325 net9531 vdd vss short_tile
xi2352 net9748 net9535 net9746 net9741 net9742 net9743 net9534 net9747 vdd vss short_tile
xi2401 net9958 net9745 net9959 net9955 net9956 net9953 net9744 net9957 vdd vss short_tile
xi2599 vdd vss enable<49> net10341 net10342 enable_tile
xi2598 vdd vss enable<48> net10304 net10305 enable_tile
xi2597 vdd vss enable<47> net10300 net10301 enable_tile
xi2596 vdd vss enable<46> net10310 net10311 enable_tile
xi2595 vdd vss enable<45> net10308 net10320 enable_tile
xi2594 vdd vss enable<44> net10315 net10316 enable_tile
xi2593 vdd vss enable<43> net10324 net10325 enable_tile
xi2592 vdd vss enable<42> net10322 net10323 enable_tile
xi2591 vdd vss enable<41> net10328 net10329 enable_tile
xi2590 vdd vss enable<40> net10337 net10338 enable_tile
xi2589 vdd vss enable<39> net10334 net10335 enable_tile
xi2588 vdd vss enable<38> net10340 net10264 enable_tile
xi2587 vdd vss enable<37> net10259 net10260 enable_tile
xi2586 vdd vss enable<36> net10269 net10270 enable_tile
xi2585 vdd vss enable<35> net10267 net10268 enable_tile
xi2584 vdd vss enable<34> net10273 net10274 enable_tile
xi2583 vdd vss enable<33> net10282 net10283 enable_tile
xi2582 vdd vss enable<32> net10279 net10280 enable_tile
xi2581 vdd vss enable<31> net10287 net10288 enable_tile
xi2580 vdd vss enable<30> net10285 net10296 enable_tile
xi2579 vdd vss enable<29> net10292 net10293 enable_tile
xi2578 vdd vss enable<28> net10297 net10298 enable_tile
xi2577 vdd vss enable<27> net10218 net10219 enable_tile
xi2576 vdd vss enable<26> net10228 net10229 enable_tile
xi2575 vdd vss enable<25> net10225 net10226 enable_tile
xi2574 vdd vss enable<24> net10233 net10234 enable_tile
xi2573 vdd vss enable<23> net10231 net10243 enable_tile
xi2572 vdd vss enable<22> net10238 net10239 enable_tile
xi2571 vdd vss enable<21> net10247 net10248 enable_tile
xi2570 vdd vss enable<20> net10245 net10246 enable_tile
xi2569 vdd vss enable<19> net10251 net10252 enable_tile
xi2568 vdd vss enable<18> net10256 net10257 enable_tile
xi2567 vdd vss enable<17> net10180 net10181 enable_tile
xi2566 vdd vss enable<16> net10178 net10190 enable_tile
xi2565 vdd vss enable<15> net10185 net10186 enable_tile
xi2564 vdd vss enable<14> net10194 net10195 enable_tile
xi2563 vdd vss enable<13> net10192 net10193 enable_tile
xi2562 vdd vss enable<12> net10198 net10199 enable_tile
xi2561 vdd vss enable<11> net10207 net10208 enable_tile
xi2560 vdd vss enable<10> net10204 net10205 enable_tile
xi2559 vdd vss enable<9> net10212 net10213 enable_tile
xi2558 vdd vss enable<8> net10210 net10216 enable_tile
xi2557 vdd vss enable<7> net10141 net10142 enable_tile
xi2556 vdd vss enable<6> net10138 net10139 enable_tile
xi2555 vdd vss enable<5> net10146 net10147 enable_tile
xi2554 vdd vss enable<4> net10155 net10156 enable_tile
xi2553 vdd vss enable<3> net10152 net10153 enable_tile
xi2552 vdd vss enable<2> net10160 net10161 enable_tile
xi2551 vdd vss enable<1> net10158 net10164 enable_tile
xi2550 vdd vss enable<0> net10167 net10168 enable_tile
xi2549 vdd vss enable<0> net10170 net10169 enable_tile
xi2548 vdd vss enable<1> net9966 net9965 enable_tile
xi2547 vdd vss enable<2> net9755 net9754 enable_tile
xi2546 vdd vss enable<3> net9551 net9550 enable_tile
xi2545 vdd vss enable<4> net9340 net9339 enable_tile
xi2544 vdd vss enable<5> net9130 net9129 enable_tile
xi2543 vdd vss enable<6> net8926 net8925 enable_tile
xi2542 vdd vss enable<7> net8716 net8715 enable_tile
xi2541 vdd vss enable<8> net8584 net8583 enable_tile
xi2540 vdd vss enable<9> net8379 net8378 enable_tile
xi2539 vdd vss enable<10> net8175 net8174 enable_tile
xi2538 vdd vss enable<11> net7964 net7963 enable_tile
xi2537 vdd vss enable<12> net7754 net7753 enable_tile
xi2536 vdd vss enable<13> net7550 net7549 enable_tile
xi2535 vdd vss enable<14> net7340 net7339 enable_tile
xi2534 vdd vss enable<15> net7129 net7128 enable_tile
xi2533 vdd vss enable<16> net6926 net6925 enable_tile
xi2532 vdd vss enable<17> net6715 net6714 enable_tile
xi2531 vdd vss enable<18> net6511 net6510 enable_tile
xi2530 vdd vss enable<19> net6379 net6378 enable_tile
xi2529 vdd vss enable<20> net6175 net6174 enable_tile
xi2528 vdd vss enable<21> net5965 net5964 enable_tile
xi2527 vdd vss enable<22> net5754 net5753 enable_tile
xi2526 vdd vss enable<23> net5551 net5550 enable_tile
xi2525 vdd vss enable<24> net5340 net5339 enable_tile
xi2524 vdd vss enable<25> net5136 net5135 enable_tile
xi2523 vdd vss enable<26> net4925 net4924 enable_tile
xi2522 vdd vss enable<27> net4712 net4713 enable_tile
xi2521 vdd vss enable<28> net4505 net4506 enable_tile
xi2520 vdd vss enable<29> net4377 net4378 enable_tile
xi2519 vdd vss enable<30> net4171 net4172 enable_tile
xi2518 vdd vss enable<31> net3962 net3963 enable_tile
xi2517 vdd vss enable<32> net3756 net3757 enable_tile
xi2516 vdd vss enable<33> net3546 net3547 enable_tile
xi2515 vdd vss enable<34> net3338 net3339 enable_tile
xi2514 vdd vss enable<35> net3132 net3133 enable_tile
xi2513 vdd vss enable<36> net1089 net1090 enable_tile
xi2512 vdd vss enable<37> net1836 net1837 enable_tile
xi2511 vdd vss enable<38> net1650 net1651 enable_tile
xi2510 vdd vss enable<39> net1951 net1952 enable_tile
xi2509 vdd vss enable<40> net2149 net2150 enable_tile
xi2508 vdd vss enable<41> net2349 net2350 enable_tile
xi2507 vdd vss enable<42> net2550 net2551 enable_tile
xi2506 vdd vss enable<43> net2749 net2750 enable_tile
xi2505 vdd vss enable<44> net2950 net2949 enable_tile
xi2504 vdd vss enable<45> net3067 net3066 enable_tile
xi2503 vdd vss enable<46> net700 net699 enable_tile
xi2502 vdd vss enable<47> net322 net321 enable_tile
xi2501 vdd vss enable<48> net1343 net1344 enable_tile
xi2500 vdd vss enable<49> net1258 net1257 enable_tile
.END
