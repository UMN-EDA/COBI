module decoder 
  (
   input wire 						    address_enable,
   input wire [$clog2(`ARRAY_SIZE)-1:0] WL_num,
   input                                prechargeb,
   output [`ARRAY_SIZE-1:0]			    WL
   );
	reg [`ARRAY_SIZE-1:0] WWL_temp;
	assign WL = WWL_temp;
	

    always @(*) begin
        if (address_enable && prechargeb) begin
            case (WL_num+1)
                 1: WWL_temp = 50'b00000000000000000000000000000000000000000000000001;
                 2: WWL_temp = 50'b00000000000000000000000000000000000000000000000010;
                 3: WWL_temp = 50'b00000000000000000000000000000000000000000000000100;
                 4: WWL_temp = 50'b00000000000000000000000000000000000000000000001000;
                 5: WWL_temp = 50'b00000000000000000000000000000000000000000000010000;
                 6: WWL_temp = 50'b00000000000000000000000000000000000000000000100000;
                 7: WWL_temp = 50'b00000000000000000000000000000000000000000001000000;
                 8: WWL_temp = 50'b00000000000000000000000000000000000000000010000000;
                 9: WWL_temp = 50'b00000000000000000000000000000000000000000100000000;
                10: WWL_temp = 50'b00000000000000000000000000000000000000001000000000;
                11: WWL_temp = 50'b00000000000000000000000000000000000000010000000000;
                12: WWL_temp = 50'b00000000000000000000000000000000000000100000000000;
                13: WWL_temp = 50'b00000000000000000000000000000000000001000000000000;
                14: WWL_temp = 50'b00000000000000000000000000000000000010000000000000;
                15: WWL_temp = 50'b00000000000000000000000000000000000100000000000000;
                16: WWL_temp = 50'b00000000000000000000000000000000001000000000000000;
                17: WWL_temp = 50'b00000000000000000000000000000000010000000000000000;
                18: WWL_temp = 50'b00000000000000000000000000000000100000000000000000;
                19: WWL_temp = 50'b00000000000000000000000000000001000000000000000000;
                20: WWL_temp = 50'b00000000000000000000000000000010000000000000000000;
                21: WWL_temp = 50'b00000000000000000000000000000100000000000000000000;
                22: WWL_temp = 50'b00000000000000000000000000001000000000000000000000;
                23: WWL_temp = 50'b00000000000000000000000000010000000000000000000000;
                24: WWL_temp = 50'b00000000000000000000000000100000000000000000000000;
                25: WWL_temp = 50'b00000000000000000000000001000000000000000000000000;
                26: WWL_temp = 50'b00000000000000000000000010000000000000000000000000;
                27: WWL_temp = 50'b00000000000000000000000100000000000000000000000000;
                28: WWL_temp = 50'b00000000000000000000001000000000000000000000000000;
                29: WWL_temp = 50'b00000000000000000000010000000000000000000000000000;
                30: WWL_temp = 50'b00000000000000000000100000000000000000000000000000;
                31: WWL_temp = 50'b00000000000000000001000000000000000000000000000000;
                32: WWL_temp = 50'b00000000000000000010000000000000000000000000000000;
                33: WWL_temp = 50'b00000000000000000100000000000000000000000000000000;
                34: WWL_temp = 50'b00000000000000001000000000000000000000000000000000;
                35: WWL_temp = 50'b00000000000000010000000000000000000000000000000000;
                36: WWL_temp = 50'b00000000000000100000000000000000000000000000000000;
                37: WWL_temp = 50'b00000000000001000000000000000000000000000000000000;
                38: WWL_temp = 50'b00000000000010000000000000000000000000000000000000;
                39: WWL_temp = 50'b00000000000100000000000000000000000000000000000000;
		        40: WWL_temp = 50'b00000000001000000000000000000000000000000000000000;
		        41: WWL_temp = 50'b00000000010000000000000000000000000000000000000000;
		        42: WWL_temp = 50'b00000000100000000000000000000000000000000000000000;
		        43: WWL_temp = 50'b00000001000000000000000000000000000000000000000000;
		        44: WWL_temp = 50'b00000010000000000000000000000000000000000000000000;
		        45: WWL_temp = 50'b00000100000000000000000000000000000000000000000000;
		        46: WWL_temp = 50'b00001000000000000000000000000000000000000000000000;
		        47: WWL_temp = 50'b00010000000000000000000000000000000000000000000000;
		        48: WWL_temp = 50'b00100000000000000000000000000000000000000000000000;
		        49: WWL_temp = 50'b01000000000000000000000000000000000000000000000000;
		        50: WWL_temp = 50'b10000000000000000000000000000000000000000000000000;
                default: WWL_temp = 50'b00000000000000000000000000000000000000000000000000;
            endcase
        end else begin
                WWL_temp = 50'b00000000000000000000000000000000000000000000000000;
        end
	end
endmodule
