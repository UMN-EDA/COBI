// define
//`define CORE 0
// AXI interface
`define DATA_WIDTH_IN_STREAM 16
`define DATA_WIDTH_OUT_STREAM 1
`define DATA_WIDTH 16
`define FIFO_IN_REG 1
`define FIFO_OUT_REG 1
`define FIFO_DEPTH 4
`define FIFO_LOG2_DEPTH 2
`define FIFO_CMD_LENGTH_IN 17
`define FIFO_CMD_LENGTH_OUT 2
`define WORD_WIDTH 4
`define SHIL 25

// axi and core
`define OUTPUT_REG_SIZE 69
`define OUTPUT_RESULT_SIZE 69
`define NUM_CONTROL 13

// Ising core
`define ARRAY_SIZE 50
`define CORE_SIZE 50



// parameter
`define M_COUNT 1
`define TOTAL_ARRAY_NUM_BIT 200 // Array_size * 4

// accelerator
`define NUM_ROW 46
`define ENERGY_WIDTH 15
`define GREDIENT_SUM_WIDTH 11
`define FAILS_WIDTH 15


